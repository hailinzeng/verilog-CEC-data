module c1355
( id_1gat ,id_8gat ,id_15gat ,id_22gat ,id_29gat ,id_36gat ,id_43gat ,id_50gat ,id_57gat ,id_64gat ,id_71gat ,id_78gat ,id_85gat ,id_92gat ,id_99gat ,id_106gat ,id_113gat ,id_120gat ,id_127gat ,id_134gat ,id_141gat ,id_148gat ,id_155gat ,id_162gat ,id_169gat ,id_176gat ,id_183gat ,id_190gat ,id_197gat ,id_204gat ,id_211gat ,id_218gat ,id_225gat ,id_226gat ,id_227gat ,id_228gat ,id_229gat ,id_230gat ,id_231gat ,id_232gat ,id_233gat ,id_1324gat ,id_1325gat ,id_1326gat ,id_1327gat ,id_1328gat ,id_1329gat ,id_1330gat ,id_1331gat ,id_1332gat ,id_1333gat ,id_1334gat ,id_1335gat ,id_1336gat ,id_1337gat ,id_1338gat ,id_1339gat ,id_1340gat ,id_1341gat ,id_1342gat ,id_1343gat ,id_1344gat ,id_1345gat ,id_1346gat ,id_1347gat ,id_1348gat ,id_1349gat ,id_1350gat ,id_1351gat ,id_1352gat ,id_1353gat ,id_1354gat ,id_1355gat );

input id_1gat, id_8gat, id_15gat, id_22gat, id_29gat, id_36gat, id_43gat, id_50gat, id_57gat, id_64gat, id_71gat, id_78gat, id_85gat, id_92gat, id_99gat, id_106gat, id_113gat, id_120gat, id_127gat, id_134gat, id_141gat, id_148gat, id_155gat, id_162gat, id_169gat, id_176gat, id_183gat, id_190gat, id_197gat, id_204gat, id_211gat, id_218gat, id_225gat, id_226gat, id_227gat, id_228gat, id_229gat, id_230gat, id_231gat, id_232gat, id_233gat;

output id_1324gat, id_1325gat, id_1326gat, id_1327gat, id_1328gat, id_1329gat, id_1330gat, id_1331gat, id_1332gat, id_1333gat, id_1334gat, id_1335gat, id_1336gat, id_1337gat, id_1338gat, id_1339gat, id_1340gat, id_1341gat, id_1342gat, id_1343gat, id_1344gat, id_1345gat, id_1346gat, id_1347gat, id_1348gat, id_1349gat, id_1350gat, id_1351gat, id_1352gat, id_1353gat, id_1354gat, id_1355gat;

and ( id_242gat, id_225gat, id_233gat);
and ( id_245gat, id_226gat, id_233gat);
and ( id_248gat, id_227gat, id_233gat);
and ( id_251gat, id_228gat, id_233gat);
and ( id_254gat, id_229gat, id_233gat);
and ( id_257gat, id_230gat, id_233gat);
and ( id_260gat, id_231gat, id_233gat);
and ( id_263gat, id_232gat, id_233gat);
nand ( id_266gat, id_1gat, id_8gat);
nand ( id_269gat, id_15gat, id_22gat);
nand ( id_272gat, id_29gat, id_36gat);
nand ( id_275gat, id_43gat, id_50gat);
nand ( id_278gat, id_57gat, id_64gat);
nand ( id_281gat, id_71gat, id_78gat);
nand ( id_284gat, id_85gat, id_92gat);
nand ( id_287gat, id_99gat, id_106gat);
nand ( id_290gat, id_113gat, id_120gat);
nand ( id_293gat, id_127gat, id_134gat);
nand ( id_296gat, id_141gat, id_148gat);
nand ( id_299gat, id_155gat, id_162gat);
nand ( id_302gat, id_169gat, id_176gat);
nand ( id_305gat, id_183gat, id_190gat);
nand ( id_308gat, id_197gat, id_204gat);
nand ( id_311gat, id_211gat, id_218gat);
nand ( id_314gat, id_1gat, id_29gat);
nand ( id_317gat, id_57gat, id_85gat);
nand ( id_320gat, id_8gat, id_36gat);
nand ( id_323gat, id_64gat, id_92gat);
nand ( id_326gat, id_15gat, id_43gat);
nand ( id_329gat, id_71gat, id_99gat);
nand ( id_332gat, id_22gat, id_50gat);
nand ( id_335gat, id_78gat, id_106gat);
nand ( id_338gat, id_113gat, id_141gat);
nand ( id_341gat, id_169gat, id_197gat);
nand ( id_344gat, id_120gat, id_148gat);
nand ( id_347gat, id_176gat, id_204gat);
nand ( id_350gat, id_127gat, id_155gat);
nand ( id_353gat, id_183gat, id_211gat);
nand ( id_356gat, id_134gat, id_162gat);
nand ( id_359gat, id_190gat, id_218gat);
nand ( id_362gat, id_1gat, id_266gat);
nand ( id_363gat, id_8gat, id_266gat);
nand ( id_364gat, id_15gat, id_269gat);
nand ( id_365gat, id_22gat, id_269gat);
nand ( id_366gat, id_29gat, id_272gat);
nand ( id_367gat, id_36gat, id_272gat);
nand ( id_368gat, id_43gat, id_275gat);
nand ( id_369gat, id_50gat, id_275gat);
nand ( id_370gat, id_57gat, id_278gat);
nand ( id_371gat, id_64gat, id_278gat);
nand ( id_372gat, id_71gat, id_281gat);
nand ( id_373gat, id_78gat, id_281gat);
nand ( id_374gat, id_85gat, id_284gat);
nand ( id_375gat, id_92gat, id_284gat);
nand ( id_376gat, id_99gat, id_287gat);
nand ( id_377gat, id_106gat, id_287gat);
nand ( id_378gat, id_113gat, id_290gat);
nand ( id_379gat, id_120gat, id_290gat);
nand ( id_380gat, id_127gat, id_293gat);
nand ( id_381gat, id_134gat, id_293gat);
nand ( id_382gat, id_141gat, id_296gat);
nand ( id_383gat, id_148gat, id_296gat);
nand ( id_384gat, id_155gat, id_299gat);
nand ( id_385gat, id_162gat, id_299gat);
nand ( id_386gat, id_169gat, id_302gat);
nand ( id_387gat, id_176gat, id_302gat);
nand ( id_388gat, id_183gat, id_305gat);
nand ( id_389gat, id_190gat, id_305gat);
nand ( id_390gat, id_197gat, id_308gat);
nand ( id_391gat, id_204gat, id_308gat);
nand ( id_392gat, id_211gat, id_311gat);
nand ( id_393gat, id_218gat, id_311gat);
nand ( id_394gat, id_1gat, id_314gat);
nand ( id_395gat, id_29gat, id_314gat);
nand ( id_396gat, id_57gat, id_317gat);
nand ( id_397gat, id_85gat, id_317gat);
nand ( id_398gat, id_8gat, id_320gat);
nand ( id_399gat, id_36gat, id_320gat);
nand ( id_400gat, id_64gat, id_323gat);
nand ( id_401gat, id_92gat, id_323gat);
nand ( id_402gat, id_15gat, id_326gat);
nand ( id_403gat, id_43gat, id_326gat);
nand ( id_404gat, id_71gat, id_329gat);
nand ( id_405gat, id_99gat, id_329gat);
nand ( id_406gat, id_22gat, id_332gat);
nand ( id_407gat, id_50gat, id_332gat);
nand ( id_408gat, id_78gat, id_335gat);
nand ( id_409gat, id_106gat, id_335gat);
nand ( id_410gat, id_113gat, id_338gat);
nand ( id_411gat, id_141gat, id_338gat);
nand ( id_412gat, id_169gat, id_341gat);
nand ( id_413gat, id_197gat, id_341gat);
nand ( id_414gat, id_120gat, id_344gat);
nand ( id_415gat, id_148gat, id_344gat);
nand ( id_416gat, id_176gat, id_347gat);
nand ( id_417gat, id_204gat, id_347gat);
nand ( id_418gat, id_127gat, id_350gat);
nand ( id_419gat, id_155gat, id_350gat);
nand ( id_420gat, id_183gat, id_353gat);
nand ( id_421gat, id_211gat, id_353gat);
nand ( id_422gat, id_134gat, id_356gat);
nand ( id_423gat, id_162gat, id_356gat);
nand ( id_424gat, id_190gat, id_359gat);
nand ( id_425gat, id_218gat, id_359gat);
nand ( id_426gat, id_362gat, id_363gat);
nand ( id_429gat, id_364gat, id_365gat);
nand ( id_432gat, id_366gat, id_367gat);
nand ( id_435gat, id_368gat, id_369gat);
nand ( id_438gat, id_370gat, id_371gat);
nand ( id_441gat, id_372gat, id_373gat);
nand ( id_444gat, id_374gat, id_375gat);
nand ( id_447gat, id_376gat, id_377gat);
nand ( id_450gat, id_378gat, id_379gat);
nand ( id_453gat, id_380gat, id_381gat);
nand ( id_456gat, id_382gat, id_383gat);
nand ( id_459gat, id_384gat, id_385gat);
nand ( id_462gat, id_386gat, id_387gat);
nand ( id_465gat, id_388gat, id_389gat);
nand ( id_468gat, id_390gat, id_391gat);
nand ( id_471gat, id_392gat, id_393gat);
nand ( id_474gat, id_394gat, id_395gat);
nand ( id_477gat, id_396gat, id_397gat);
nand ( id_480gat, id_398gat, id_399gat);
nand ( id_483gat, id_400gat, id_401gat);
nand ( id_486gat, id_402gat, id_403gat);
nand ( id_489gat, id_404gat, id_405gat);
nand ( id_492gat, id_406gat, id_407gat);
nand ( id_495gat, id_408gat, id_409gat);
nand ( id_498gat, id_410gat, id_411gat);
nand ( id_501gat, id_412gat, id_413gat);
nand ( id_504gat, id_414gat, id_415gat);
nand ( id_507gat, id_416gat, id_417gat);
nand ( id_510gat, id_418gat, id_419gat);
nand ( id_513gat, id_420gat, id_421gat);
nand ( id_516gat, id_422gat, id_423gat);
nand ( id_519gat, id_424gat, id_425gat);
nand ( id_522gat, id_426gat, id_429gat);
nand ( id_525gat, id_432gat, id_435gat);
nand ( id_528gat, id_438gat, id_441gat);
nand ( id_531gat, id_444gat, id_447gat);
nand ( id_534gat, id_450gat, id_453gat);
nand ( id_537gat, id_456gat, id_459gat);
nand ( id_540gat, id_462gat, id_465gat);
nand ( id_543gat, id_468gat, id_471gat);
nand ( id_546gat, id_474gat, id_477gat);
nand ( id_549gat, id_480gat, id_483gat);
nand ( id_552gat, id_486gat, id_489gat);
nand ( id_555gat, id_492gat, id_495gat);
nand ( id_558gat, id_498gat, id_501gat);
nand ( id_561gat, id_504gat, id_507gat);
nand ( id_564gat, id_510gat, id_513gat);
nand ( id_567gat, id_516gat, id_519gat);
nand ( id_570gat, id_426gat, id_522gat);
nand ( id_571gat, id_429gat, id_522gat);
nand ( id_572gat, id_432gat, id_525gat);
nand ( id_573gat, id_435gat, id_525gat);
nand ( id_574gat, id_438gat, id_528gat);
nand ( id_575gat, id_441gat, id_528gat);
nand ( id_576gat, id_444gat, id_531gat);
nand ( id_577gat, id_447gat, id_531gat);
nand ( id_578gat, id_450gat, id_534gat);
nand ( id_579gat, id_453gat, id_534gat);
nand ( id_580gat, id_456gat, id_537gat);
nand ( id_581gat, id_459gat, id_537gat);
nand ( id_582gat, id_462gat, id_540gat);
nand ( id_583gat, id_465gat, id_540gat);
nand ( id_584gat, id_468gat, id_543gat);
nand ( id_585gat, id_471gat, id_543gat);
nand ( id_586gat, id_474gat, id_546gat);
nand ( id_587gat, id_477gat, id_546gat);
nand ( id_588gat, id_480gat, id_549gat);
nand ( id_589gat, id_483gat, id_549gat);
nand ( id_590gat, id_486gat, id_552gat);
nand ( id_591gat, id_489gat, id_552gat);
nand ( id_592gat, id_492gat, id_555gat);
nand ( id_593gat, id_495gat, id_555gat);
nand ( id_594gat, id_498gat, id_558gat);
nand ( id_595gat, id_501gat, id_558gat);
nand ( id_596gat, id_504gat, id_561gat);
nand ( id_597gat, id_507gat, id_561gat);
nand ( id_598gat, id_510gat, id_564gat);
nand ( id_599gat, id_513gat, id_564gat);
nand ( id_600gat, id_516gat, id_567gat);
nand ( id_601gat, id_519gat, id_567gat);
nand ( id_602gat, id_570gat, id_571gat);
nand ( id_607gat, id_572gat, id_573gat);
nand ( id_612gat, id_574gat, id_575gat);
nand ( id_617gat, id_576gat, id_577gat);
nand ( id_622gat, id_578gat, id_579gat);
nand ( id_627gat, id_580gat, id_581gat);
nand ( id_632gat, id_582gat, id_583gat);
nand ( id_637gat, id_584gat, id_585gat);
nand ( id_642gat, id_586gat, id_587gat);
nand ( id_645gat, id_588gat, id_589gat);
nand ( id_648gat, id_590gat, id_591gat);
nand ( id_651gat, id_592gat, id_593gat);
nand ( id_654gat, id_594gat, id_595gat);
nand ( id_657gat, id_596gat, id_597gat);
nand ( id_660gat, id_598gat, id_599gat);
nand ( id_663gat, id_600gat, id_601gat);
nand ( id_666gat, id_602gat, id_607gat);
nand ( id_669gat, id_612gat, id_617gat);
nand ( id_672gat, id_602gat, id_612gat);
nand ( id_675gat, id_607gat, id_617gat);
nand ( id_678gat, id_622gat, id_627gat);
nand ( id_681gat, id_632gat, id_637gat);
nand ( id_684gat, id_622gat, id_632gat);
nand ( id_687gat, id_627gat, id_637gat);
nand ( id_690gat, id_602gat, id_666gat);
nand ( id_691gat, id_607gat, id_666gat);
nand ( id_692gat, id_612gat, id_669gat);
nand ( id_693gat, id_617gat, id_669gat);
nand ( id_694gat, id_602gat, id_672gat);
nand ( id_695gat, id_612gat, id_672gat);
nand ( id_696gat, id_607gat, id_675gat);
nand ( id_697gat, id_617gat, id_675gat);
nand ( id_698gat, id_622gat, id_678gat);
nand ( id_699gat, id_627gat, id_678gat);
nand ( id_700gat, id_632gat, id_681gat);
nand ( id_701gat, id_637gat, id_681gat);
nand ( id_702gat, id_622gat, id_684gat);
nand ( id_703gat, id_632gat, id_684gat);
nand ( id_704gat, id_627gat, id_687gat);
nand ( id_705gat, id_637gat, id_687gat);
nand ( id_706gat, id_690gat, id_691gat);
nand ( id_709gat, id_692gat, id_693gat);
nand ( id_712gat, id_694gat, id_695gat);
nand ( id_715gat, id_696gat, id_697gat);
nand ( id_718gat, id_698gat, id_699gat);
nand ( id_721gat, id_700gat, id_701gat);
nand ( id_724gat, id_702gat, id_703gat);
nand ( id_727gat, id_704gat, id_705gat);
nand ( id_730gat, id_242gat, id_718gat);
nand ( id_733gat, id_245gat, id_721gat);
nand ( id_736gat, id_248gat, id_724gat);
nand ( id_739gat, id_251gat, id_727gat);
nand ( id_742gat, id_254gat, id_706gat);
nand ( id_745gat, id_257gat, id_709gat);
nand ( id_748gat, id_260gat, id_712gat);
nand ( id_751gat, id_263gat, id_715gat);
nand ( id_754gat, id_242gat, id_730gat);
nand ( id_755gat, id_718gat, id_730gat);
nand ( id_756gat, id_245gat, id_733gat);
nand ( id_757gat, id_721gat, id_733gat);
nand ( id_758gat, id_248gat, id_736gat);
nand ( id_759gat, id_724gat, id_736gat);
nand ( id_760gat, id_251gat, id_739gat);
nand ( id_761gat, id_727gat, id_739gat);
nand ( id_762gat, id_254gat, id_742gat);
nand ( id_763gat, id_706gat, id_742gat);
nand ( id_764gat, id_257gat, id_745gat);
nand ( id_765gat, id_709gat, id_745gat);
nand ( id_766gat, id_260gat, id_748gat);
nand ( id_767gat, id_712gat, id_748gat);
nand ( id_768gat, id_263gat, id_751gat);
nand ( id_769gat, id_715gat, id_751gat);
nand ( id_770gat, id_754gat, id_755gat);
nand ( id_773gat, id_756gat, id_757gat);
nand ( id_776gat, id_758gat, id_759gat);
nand ( id_779gat, id_760gat, id_761gat);
nand ( id_782gat, id_762gat, id_763gat);
nand ( id_785gat, id_764gat, id_765gat);
nand ( id_788gat, id_766gat, id_767gat);
nand ( id_791gat, id_768gat, id_769gat);
nand ( id_794gat, id_642gat, id_770gat);
nand ( id_797gat, id_645gat, id_773gat);
nand ( id_800gat, id_648gat, id_776gat);
nand ( id_803gat, id_651gat, id_779gat);
nand ( id_806gat, id_654gat, id_782gat);
nand ( id_809gat, id_657gat, id_785gat);
nand ( id_812gat, id_660gat, id_788gat);
nand ( id_815gat, id_663gat, id_791gat);
nand ( id_818gat, id_642gat, id_794gat);
nand ( id_819gat, id_770gat, id_794gat);
nand ( id_820gat, id_645gat, id_797gat);
nand ( id_821gat, id_773gat, id_797gat);
nand ( id_822gat, id_648gat, id_800gat);
nand ( id_823gat, id_776gat, id_800gat);
nand ( id_824gat, id_651gat, id_803gat);
nand ( id_825gat, id_779gat, id_803gat);
nand ( id_826gat, id_654gat, id_806gat);
nand ( id_827gat, id_782gat, id_806gat);
nand ( id_828gat, id_657gat, id_809gat);
nand ( id_829gat, id_785gat, id_809gat);
nand ( id_830gat, id_660gat, id_812gat);
nand ( id_831gat, id_788gat, id_812gat);
nand ( id_832gat, id_663gat, id_815gat);
nand ( id_833gat, id_791gat, id_815gat);
nand ( id_834gat, id_818gat, id_819gat);
nand ( id_847gat, id_820gat, id_821gat);
nand ( id_860gat, id_822gat, id_823gat);
nand ( id_873gat, id_824gat, id_825gat);
nand ( id_886gat, id_828gat, id_829gat);
nand ( id_899gat, id_832gat, id_833gat);
nand ( id_912gat, id_830gat, id_831gat);
nand ( id_925gat, id_826gat, id_827gat);
not ( id_938gat, id_834gat);
not ( id_939gat, id_847gat);
not ( id_940gat, id_860gat);
not ( id_941gat, id_834gat);
not ( id_942gat, id_847gat);
not ( id_943gat, id_873gat);
not ( id_944gat, id_834gat);
not ( id_945gat, id_860gat);
not ( id_946gat, id_873gat);
not ( id_947gat, id_847gat);
not ( id_948gat, id_860gat);
not ( id_949gat, id_873gat);
not ( id_950gat, id_886gat);
not ( id_951gat, id_899gat);
not ( id_952gat, id_886gat);
not ( id_953gat, id_912gat);
not ( id_954gat, id_925gat);
not ( id_955gat, id_899gat);
not ( id_956gat, id_925gat);
not ( id_957gat, id_912gat);
not ( id_958gat, id_925gat);
not ( id_959gat, id_886gat);
not ( id_960gat, id_912gat);
not ( id_961gat, id_925gat);
not ( id_962gat, id_886gat);
not ( id_963gat, id_899gat);
not ( id_964gat, id_925gat);
not ( id_965gat, id_912gat);
not ( id_966gat, id_899gat);
not ( id_967gat, id_886gat);
not ( id_968gat, id_912gat);
not ( id_969gat, id_899gat);
not ( id_970gat, id_847gat);
not ( id_971gat, id_873gat);
not ( id_972gat, id_847gat);
not ( id_973gat, id_860gat);
not ( id_974gat, id_834gat);
not ( id_975gat, id_873gat);
not ( id_976gat, id_834gat);
not ( id_977gat, id_860gat);
and ( id_978gat, id_938gat, id_939gat, id_940gat, id_873gat);
and ( id_979gat, id_941gat, id_942gat, id_860gat, id_943gat);
and ( id_980gat, id_944gat, id_847gat, id_945gat, id_946gat);
and ( id_981gat, id_834gat, id_947gat, id_948gat, id_949gat);
and ( id_982gat, id_958gat, id_959gat, id_960gat, id_899gat);
and ( id_983gat, id_961gat, id_962gat, id_912gat, id_963gat);
and ( id_984gat, id_964gat, id_886gat, id_965gat, id_966gat);
and ( id_985gat, id_925gat, id_967gat, id_968gat, id_969gat);
or ( id_986gat, id_978gat, id_979gat, id_980gat, id_981gat);
or ( id_991gat, id_982gat, id_983gat, id_984gat, id_985gat);
and ( id_996gat, id_925gat, id_950gat, id_912gat, id_951gat, id_986gat);
and ( id_1001gat, id_925gat, id_952gat, id_953gat, id_899gat, id_986gat);
and ( id_1006gat, id_954gat, id_886gat, id_912gat, id_955gat, id_986gat);
and ( id_1011gat, id_956gat, id_886gat, id_957gat, id_899gat, id_986gat);
and ( id_1016gat, id_834gat, id_970gat, id_860gat, id_971gat, id_991gat);
and ( id_1021gat, id_834gat, id_972gat, id_973gat, id_873gat, id_991gat);
and ( id_1026gat, id_974gat, id_847gat, id_860gat, id_975gat, id_991gat);
and ( id_1031gat, id_976gat, id_847gat, id_977gat, id_873gat, id_991gat);
and ( id_1036gat, id_834gat, id_996gat);
and ( id_1039gat, id_847gat, id_996gat);
and ( id_1042gat, id_860gat, id_996gat);
and ( id_1045gat, id_873gat, id_996gat);
and ( id_1048gat, id_834gat, id_1001gat);
and ( id_1051gat, id_847gat, id_1001gat);
and ( id_1054gat, id_860gat, id_1001gat);
and ( id_1057gat, id_873gat, id_1001gat);
and ( id_1060gat, id_834gat, id_1006gat);
and ( id_1063gat, id_847gat, id_1006gat);
and ( id_1066gat, id_860gat, id_1006gat);
and ( id_1069gat, id_873gat, id_1006gat);
and ( id_1072gat, id_834gat, id_1011gat);
and ( id_1075gat, id_847gat, id_1011gat);
and ( id_1078gat, id_860gat, id_1011gat);
and ( id_1081gat, id_873gat, id_1011gat);
and ( id_1084gat, id_925gat, id_1016gat);
and ( id_1087gat, id_886gat, id_1016gat);
and ( id_1090gat, id_912gat, id_1016gat);
and ( id_1093gat, id_899gat, id_1016gat);
and ( id_1096gat, id_925gat, id_1021gat);
and ( id_1099gat, id_886gat, id_1021gat);
and ( id_1102gat, id_912gat, id_1021gat);
and ( id_1105gat, id_899gat, id_1021gat);
and ( id_1108gat, id_925gat, id_1026gat);
and ( id_1111gat, id_886gat, id_1026gat);
and ( id_1114gat, id_912gat, id_1026gat);
and ( id_1117gat, id_899gat, id_1026gat);
and ( id_1120gat, id_925gat, id_1031gat);
and ( id_1123gat, id_886gat, id_1031gat);
and ( id_1126gat, id_912gat, id_1031gat);
and ( id_1129gat, id_899gat, id_1031gat);
nand ( id_1132gat, id_1gat, id_1036gat);
nand ( id_1135gat, id_8gat, id_1039gat);
nand ( id_1138gat, id_15gat, id_1042gat);
nand ( id_1141gat, id_22gat, id_1045gat);
nand ( id_1144gat, id_29gat, id_1048gat);
nand ( id_1147gat, id_36gat, id_1051gat);
nand ( id_1150gat, id_43gat, id_1054gat);
nand ( id_1153gat, id_50gat, id_1057gat);
nand ( id_1156gat, id_57gat, id_1060gat);
nand ( id_1159gat, id_64gat, id_1063gat);
nand ( id_1162gat, id_71gat, id_1066gat);
nand ( id_1165gat, id_78gat, id_1069gat);
nand ( id_1168gat, id_85gat, id_1072gat);
nand ( id_1171gat, id_92gat, id_1075gat);
nand ( id_1174gat, id_99gat, id_1078gat);
nand ( id_1177gat, id_106gat, id_1081gat);
nand ( id_1180gat, id_113gat, id_1084gat);
nand ( id_1183gat, id_120gat, id_1087gat);
nand ( id_1186gat, id_127gat, id_1090gat);
nand ( id_1189gat, id_134gat, id_1093gat);
nand ( id_1192gat, id_141gat, id_1096gat);
nand ( id_1195gat, id_148gat, id_1099gat);
nand ( id_1198gat, id_155gat, id_1102gat);
nand ( id_1201gat, id_162gat, id_1105gat);
nand ( id_1204gat, id_169gat, id_1108gat);
nand ( id_1207gat, id_176gat, id_1111gat);
nand ( id_1210gat, id_183gat, id_1114gat);
nand ( id_1213gat, id_190gat, id_1117gat);
nand ( id_1216gat, id_197gat, id_1120gat);
nand ( id_1219gat, id_204gat, id_1123gat);
nand ( id_1222gat, id_211gat, id_1126gat);
nand ( id_1225gat, id_218gat, id_1129gat);
nand ( id_1228gat, id_1gat, id_1132gat);
nand ( id_1229gat, id_1036gat, id_1132gat);
nand ( id_1230gat, id_8gat, id_1135gat);
nand ( id_1231gat, id_1039gat, id_1135gat);
nand ( id_1232gat, id_15gat, id_1138gat);
nand ( id_1233gat, id_1042gat, id_1138gat);
nand ( id_1234gat, id_22gat, id_1141gat);
nand ( id_1235gat, id_1045gat, id_1141gat);
nand ( id_1236gat, id_29gat, id_1144gat);
nand ( id_1237gat, id_1048gat, id_1144gat);
nand ( id_1238gat, id_36gat, id_1147gat);
nand ( id_1239gat, id_1051gat, id_1147gat);
nand ( id_1240gat, id_43gat, id_1150gat);
nand ( id_1241gat, id_1054gat, id_1150gat);
nand ( id_1242gat, id_50gat, id_1153gat);
nand ( id_1243gat, id_1057gat, id_1153gat);
nand ( id_1244gat, id_57gat, id_1156gat);
nand ( id_1245gat, id_1060gat, id_1156gat);
nand ( id_1246gat, id_64gat, id_1159gat);
nand ( id_1247gat, id_1063gat, id_1159gat);
nand ( id_1248gat, id_71gat, id_1162gat);
nand ( id_1249gat, id_1066gat, id_1162gat);
nand ( id_1250gat, id_78gat, id_1165gat);
nand ( id_1251gat, id_1069gat, id_1165gat);
nand ( id_1252gat, id_85gat, id_1168gat);
nand ( id_1253gat, id_1072gat, id_1168gat);
nand ( id_1254gat, id_92gat, id_1171gat);
nand ( id_1255gat, id_1075gat, id_1171gat);
nand ( id_1256gat, id_99gat, id_1174gat);
nand ( id_1257gat, id_1078gat, id_1174gat);
nand ( id_1258gat, id_106gat, id_1177gat);
nand ( id_1259gat, id_1081gat, id_1177gat);
nand ( id_1260gat, id_113gat, id_1180gat);
nand ( id_1261gat, id_1084gat, id_1180gat);
nand ( id_1262gat, id_120gat, id_1183gat);
nand ( id_1263gat, id_1087gat, id_1183gat);
nand ( id_1264gat, id_127gat, id_1186gat);
nand ( id_1265gat, id_1090gat, id_1186gat);
nand ( id_1266gat, id_134gat, id_1189gat);
nand ( id_1267gat, id_1093gat, id_1189gat);
nand ( id_1268gat, id_141gat, id_1192gat);
nand ( id_1269gat, id_1096gat, id_1192gat);
nand ( id_1270gat, id_148gat, id_1195gat);
nand ( id_1271gat, id_1099gat, id_1195gat);
nand ( id_1272gat, id_155gat, id_1198gat);
nand ( id_1273gat, id_1102gat, id_1198gat);
nand ( id_1274gat, id_162gat, id_1201gat);
nand ( id_1275gat, id_1105gat, id_1201gat);
nand ( id_1276gat, id_169gat, id_1204gat);
nand ( id_1277gat, id_1108gat, id_1204gat);
nand ( id_1278gat, id_176gat, id_1207gat);
nand ( id_1279gat, id_1111gat, id_1207gat);
nand ( id_1280gat, id_183gat, id_1210gat);
nand ( id_1281gat, id_1114gat, id_1210gat);
nand ( id_1282gat, id_190gat, id_1213gat);
nand ( id_1283gat, id_1117gat, id_1213gat);
nand ( id_1284gat, id_197gat, id_1216gat);
nand ( id_1285gat, id_1120gat, id_1216gat);
nand ( id_1286gat, id_204gat, id_1219gat);
nand ( id_1287gat, id_1123gat, id_1219gat);
nand ( id_1288gat, id_211gat, id_1222gat);
nand ( id_1289gat, id_1126gat, id_1222gat);
nand ( id_1290gat, id_218gat, id_1225gat);
nand ( id_1291gat, id_1129gat, id_1225gat);
nand ( id_1292gat, id_1228gat, id_1229gat);
nand ( id_1293gat, id_1230gat, id_1231gat);
nand ( id_1294gat, id_1232gat, id_1233gat);
nand ( id_1295gat, id_1234gat, id_1235gat);
nand ( id_1296gat, id_1236gat, id_1237gat);
nand ( id_1297gat, id_1238gat, id_1239gat);
nand ( id_1298gat, id_1240gat, id_1241gat);
nand ( id_1299gat, id_1242gat, id_1243gat);
nand ( id_1300gat, id_1244gat, id_1245gat);
nand ( id_1301gat, id_1246gat, id_1247gat);
nand ( id_1302gat, id_1248gat, id_1249gat);
nand ( id_1303gat, id_1250gat, id_1251gat);
nand ( id_1304gat, id_1252gat, id_1253gat);
nand ( id_1305gat, id_1254gat, id_1255gat);
nand ( id_1306gat, id_1256gat, id_1257gat);
nand ( id_1307gat, id_1258gat, id_1259gat);
nand ( id_1308gat, id_1260gat, id_1261gat);
nand ( id_1309gat, id_1262gat, id_1263gat);
nand ( id_1310gat, id_1264gat, id_1265gat);
nand ( id_1311gat, id_1266gat, id_1267gat);
nand ( id_1312gat, id_1268gat, id_1269gat);
nand ( id_1313gat, id_1270gat, id_1271gat);
nand ( id_1314gat, id_1272gat, id_1273gat);
nand ( id_1315gat, id_1274gat, id_1275gat);
nand ( id_1316gat, id_1276gat, id_1277gat);
nand ( id_1317gat, id_1278gat, id_1279gat);
nand ( id_1318gat, id_1280gat, id_1281gat);
nand ( id_1319gat, id_1282gat, id_1283gat);
nand ( id_1320gat, id_1284gat, id_1285gat);
nand ( id_1321gat, id_1286gat, id_1287gat);
nand ( id_1322gat, id_1288gat, id_1289gat);
nand ( id_1323gat, id_1290gat, id_1291gat);
buf ( id_1324gat, id_1292gat);
buf ( id_1325gat, id_1293gat);
buf ( id_1326gat, id_1294gat);
buf ( id_1327gat, id_1295gat);
buf ( id_1328gat, id_1296gat);
buf ( id_1329gat, id_1297gat);
buf ( id_1330gat, id_1298gat);
buf ( id_1331gat, id_1299gat);
buf ( id_1332gat, id_1300gat);
buf ( id_1333gat, id_1301gat);
buf ( id_1334gat, id_1302gat);
buf ( id_1335gat, id_1303gat);
buf ( id_1336gat, id_1304gat);
buf ( id_1337gat, id_1305gat);
buf ( id_1338gat, id_1306gat);
buf ( id_1339gat, id_1307gat);
buf ( id_1340gat, id_1308gat);
buf ( id_1341gat, id_1309gat);
buf ( id_1342gat, id_1310gat);
buf ( id_1343gat, id_1311gat);
buf ( id_1344gat, id_1312gat);
buf ( id_1345gat, id_1313gat);
buf ( id_1346gat, id_1314gat);
buf ( id_1347gat, id_1315gat);
buf ( id_1348gat, id_1316gat);
buf ( id_1349gat, id_1317gat);
buf ( id_1350gat, id_1318gat);
buf ( id_1351gat, id_1319gat);
buf ( id_1352gat, id_1320gat);
buf ( id_1353gat, id_1321gat);
buf ( id_1354gat, id_1322gat);
buf ( id_1355gat, id_1323gat);

endmodule
