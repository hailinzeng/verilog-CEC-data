module c1908nr
( id_101 ,id_104 ,id_107 ,id_110 ,id_113 ,id_116 ,id_119 ,id_122 ,id_125 ,id_128 ,id_131 ,id_134 ,id_137 ,id_140 ,id_143 ,id_146 ,id_210 ,id_214 ,id_217 ,id_221 ,id_224 ,id_227 ,id_234 ,id_237 ,id_469 ,id_472 ,id_475 ,id_478 ,id_898 ,id_900 ,id_902 ,id_952 ,id_953 ,id_3 ,id_6 ,id_9 ,id_12 ,id_30 ,id_45 ,id_48 ,id_15 ,id_18 ,id_21 ,id_24 ,id_27 ,id_33 ,id_36 ,id_39 ,id_42 ,id_75 ,id_51 ,id_54 ,id_60 ,id_63 ,id_66 ,id_69 ,id_72 ,id_57  );

input id_101, id_104, id_107, id_110, id_113, id_116, id_119, id_122, id_125, id_128, id_131, id_134, id_137, id_140, id_143, id_146, id_210, id_214, id_217, id_221, id_224, id_227, id_234, id_237, id_469, id_472, id_475, id_478, id_898, id_900, id_902, id_952, id_953;

output id_3, id_6, id_9, id_12, id_30, id_45, id_48, id_15, id_18, id_21, id_24, id_27, id_33, id_36, id_39, id_42, id_75, id_51, id_54, id_60, id_63, id_66, id_69, id_72, id_57;

not ( id_149, id_101);
not ( id_153, id_104);
not ( id_156, id_107);
not ( id_160, id_110);
not ( id_165, id_113);
not ( id_168, id_116);
not ( id_171, id_119);
not ( id_175, id_122);
not ( id_179, id_125);
not ( id_184, id_128);
not ( id_188, id_131);
not ( id_191, id_134);
not ( id_194, id_137);
not ( id_198, id_140);
not ( id_202, id_143);
not ( id_206, id_146);
nand ( id_231, id_224, id_898);
nand ( id_233, id_227, id_900);
not ( id_241, id_237);
not ( id_244, id_237);
buf ( id_245, id_234);
buf ( id_248, id_234);
not ( id_517, id_469);
not ( id_529, id_472);
not ( id_541, id_475);
not ( id_553, id_478);
not ( id_859, id_953);
not ( id_862, id_953);
not ( id_907, id_898);
not ( id_909, id_900);
buf ( id_911, id_902);
not ( id_918, id_902);
buf ( id_919, id_902);
not ( id_922, id_902);
buf ( id_926, id_952);
not ( id_930, id_952);
not ( id_932, id_952);
buf ( id_934, id_953);
not ( id_938, id_953);
buf ( id_943, id_953);
buf ( id_947, id_953);
not ( id_949, id_953);
buf ( id_1506, id_101);
buf ( id_1514, id_104);
buf ( id_1522, id_107);
buf ( id_1530, id_110);
buf ( id_1538, id_113);
buf ( id_1546, id_116);
buf ( id_1554, id_119);
buf ( id_1562, id_122);
buf ( id_1570, id_125);
buf ( id_1578, id_128);
buf ( id_1586, id_131);
buf ( id_1594, id_134);
buf ( id_1602, id_137);
buf ( id_1610, id_140);
buf ( id_1618, id_143);
buf ( id_1626, id_146);
not ( id_1512, id_1506);
not ( id_1520, id_1514);
not ( id_1528, id_1522);
not ( id_1536, id_1530);
not ( id_1544, id_1538);
not ( id_1552, id_1546);
not ( id_1560, id_1554);
not ( id_1568, id_1562);
not ( id_1576, id_1570);
not ( id_1584, id_1578);
not ( id_1592, id_1586);
not ( id_1600, id_1594);
not ( id_1608, id_1602);
not ( id_1616, id_1610);
not ( id_1624, id_1618);
not ( id_1632, id_1626);
nand ( id_50, id_930, id_947);
nand ( id_52, id_930, id_947);
nand ( id_56, id_930, id_947);
nand ( id_58, id_930, id_947);
nand ( id_62, id_930, id_947);
nand ( id_64, id_930, id_947);
buf ( id_251, id_149);
buf ( id_254, id_153);
buf ( id_288, id_165);
buf ( id_291, id_168);
buf ( id_299, id_184);
buf ( id_302, id_202);
and ( id_318, id_224, id_938);
buf ( id_321, id_179);
buf ( id_327, id_188);
buf ( id_330, id_191);
and ( id_352, id_227, id_938);
buf ( id_355, id_198);
and ( id_369, id_210, id_241, id_938);
buf ( id_382, id_206);
buf ( id_385, id_198);
nand ( id_853, id_943, id_907);
nand ( id_856, id_943, id_909);
nand ( id_893, id_248, id_237);
nand ( id_954, id_248, id_922);
nand ( id_955, id_244, id_922);
buf ( id_1050, id_160);
buf ( id_1053, id_175);
buf ( id_1176, id_179);
buf ( id_1179, id_198);
buf ( id_1197, id_149);
buf ( id_1207, id_149);
buf ( id_1222, id_153);
buf ( id_1244, id_188);
buf ( id_1278, id_156);
and ( id_1290, id_217, id_245, id_938);
buf ( id_1300, id_191);
buf ( id_1312, id_160);
buf ( id_1332, id_194);
and ( id_1335, id_221, id_245, id_938);
buf ( id_1442, id_517);
buf ( id_1450, id_517);
buf ( id_1458, id_529);
buf ( id_1466, id_529);
buf ( id_1474, id_541);
buf ( id_1482, id_541);
buf ( id_1490, id_553);
buf ( id_1498, id_553);
and ( id_1634, id_231, id_934);
and ( id_1644, id_233, id_934);
buf ( id_1657, id_156);
buf ( id_1665, id_156);
buf ( id_1697, id_171);
buf ( id_1705, id_171);
buf ( id_1713, id_206);
buf ( id_1721, id_206);
buf ( id_1745, id_194);
buf ( id_1753, id_194);
buf ( id_1785, id_160);
buf ( id_1793, id_160);
buf ( id_1814, id_165);
buf ( id_1817, id_175);
and ( id_1830, id_214, id_241, id_938);
buf ( id_1833, id_202);
buf ( id_1841, id_179);
buf ( id_1849, id_179);
buf ( id_1854, id_168);
buf ( id_1857, id_175);
buf ( id_1870, id_184);
buf ( id_1873, id_202);
buf ( id_1878, id_171);
buf ( id_1881, id_184);
not ( id_1642, id_1634);
not ( id_1652, id_1644);
not ( id_1056, id_1050);
not ( id_1057, id_1053);
not ( id_1182, id_1176);
not ( id_1183, id_1179);
not ( id_1211, id_1207);
not ( id_1298, id_1290);
not ( id_1320, id_1312);
not ( id_1338, id_1332);
not ( id_1339, id_1335);
buf ( id_457, id_210);
buf ( id_459, id_217);
nand ( id_482, id_214, id_955);
nand ( id_487, id_221, id_954);
nand ( id_492, id_210, id_955);
nand ( id_505, id_217, id_954);
not ( id_1456, id_1450);
not ( id_1448, id_1442);
not ( id_1472, id_1466);
not ( id_1464, id_1458);
not ( id_1488, id_1482);
not ( id_1480, id_1474);
not ( id_1504, id_1498);
not ( id_1496, id_1490);
nand ( id_956, id_907, id_919, id_943, id_893);
nand ( id_967, id_909, id_919, id_943, id_893);
nand ( id_978, id_926, id_949, id_893);
buf ( id_979, id_893);
buf ( id_980, id_251);
not ( id_1661, id_1657);
buf ( id_990, id_251);
not ( id_1669, id_1665);
buf ( id_1030, id_288);
not ( id_1701, id_1697);
buf ( id_1040, id_288);
not ( id_1709, id_1705);
buf ( id_1058, id_299);
not ( id_1717, id_1713);
buf ( id_1068, id_299);
not ( id_1725, id_1721);
buf ( id_1078, id_318);
buf ( id_1090, id_318);
buf ( id_1100, id_327);
not ( id_1749, id_1745);
buf ( id_1112, id_327);
not ( id_1757, id_1753);
buf ( id_1154, id_352);
not ( id_1789, id_1785);
buf ( id_1166, id_352);
not ( id_1797, id_1793);
buf ( id_1194, id_369);
not ( id_1201, id_1197);
buf ( id_1204, id_369);
not ( id_1820, id_1814);
not ( id_1821, id_1817);
not ( id_1230, id_1222);
not ( id_1836, id_1830);
not ( id_1837, id_1833);
not ( id_1252, id_1244);
buf ( id_1256, id_382);
not ( id_1845, id_1841);
buf ( id_1268, id_382);
not ( id_1853, id_1849);
not ( id_1860, id_1854);
not ( id_1861, id_1857);
not ( id_1286, id_1278);
not ( id_1876, id_1870);
not ( id_1877, id_1873);
not ( id_1308, id_1300);
not ( id_1884, id_1878);
not ( id_1885, id_1881);
buf ( id_1654, id_254);
buf ( id_1662, id_254);
buf ( id_1694, id_291);
buf ( id_1702, id_291);
buf ( id_1710, id_302);
buf ( id_1718, id_302);
buf ( id_1726, id_321);
buf ( id_1734, id_321);
buf ( id_1742, id_330);
buf ( id_1750, id_330);
buf ( id_1782, id_355);
buf ( id_1790, id_355);
buf ( id_1838, id_385);
buf ( id_1846, id_385);
nand ( id_297, id_1053, id_1056);
nand ( id_298, id_1050, id_1057);
nand ( id_361, id_1179, id_1182);
nand ( id_362, id_1176, id_1183);
nand ( id_404, id_1335, id_1338);
nand ( id_405, id_1332, id_1339);
nand ( id_1225, id_1817, id_1820);
nand ( id_1226, id_1814, id_1821);
nand ( id_1247, id_1833, id_1836);
nand ( id_1248, id_1830, id_1837);
nand ( id_1281, id_1857, id_1860);
nand ( id_1282, id_1854, id_1861);
nand ( id_1303, id_1873, id_1876);
nand ( id_1304, id_1870, id_1877);
nand ( id_1315, id_1881, id_1884);
nand ( id_1316, id_1878, id_1885);
not ( id_998, id_990);
not ( id_988, id_980);
nand ( id_268, id_297, id_298);
not ( id_1038, id_1030);
not ( id_1048, id_1040);
not ( id_1076, id_1068);
not ( id_1066, id_1058);
not ( id_1098, id_1090);
not ( id_1120, id_1112);
not ( id_1174, id_1166);
nand ( id_363, id_361, id_362);
not ( id_1210, id_1204);
nand ( id_373, id_1204, id_1211);
not ( id_1276, id_1268);
nand ( id_406, id_404, id_405);
buf ( id_566, id_482);
buf ( id_615, id_487);
nand ( id_958, id_956, id_978);
nand ( id_969, id_967, id_978);
not ( id_1660, id_1654);
nand ( id_984, id_1654, id_1661);
not ( id_1668, id_1662);
nand ( id_994, id_1662, id_1669);
not ( id_1700, id_1694);
nand ( id_1034, id_1694, id_1701);
not ( id_1708, id_1702);
nand ( id_1044, id_1702, id_1709);
not ( id_1716, id_1710);
nand ( id_1062, id_1710, id_1717);
not ( id_1724, id_1718);
nand ( id_1072, id_1718, id_1725);
not ( id_1732, id_1726);
not ( id_1086, id_1078);
not ( id_1740, id_1734);
not ( id_1748, id_1742);
nand ( id_1104, id_1742, id_1749);
not ( id_1108, id_1100);
not ( id_1756, id_1750);
nand ( id_1116, id_1750, id_1757);
not ( id_1788, id_1782);
nand ( id_1158, id_1782, id_1789);
not ( id_1162, id_1154);
not ( id_1796, id_1790);
nand ( id_1170, id_1790, id_1797);
not ( id_1200, id_1194);
nand ( id_1203, id_1194, id_1201);
nand ( id_1227, id_1225, id_1226);
nand ( id_1249, id_1247, id_1248);
not ( id_1844, id_1838);
nand ( id_1260, id_1838, id_1845);
not ( id_1264, id_1256);
not ( id_1852, id_1846);
nand ( id_1272, id_1846, id_1853);
nand ( id_1283, id_1281, id_1282);
nand ( id_1305, id_1303, id_1304);
nand ( id_1317, id_1315, id_1316);
buf ( id_1410, id_492);
buf ( id_1418, id_492);
buf ( id_1426, id_505);
buf ( id_1434, id_505);
not ( id_269, id_268);
nand ( id_372, id_1207, id_1210);
nand ( id_983, id_1657, id_1660);
nand ( id_993, id_1665, id_1668);
nand ( id_1033, id_1697, id_1700);
nand ( id_1043, id_1705, id_1708);
nand ( id_1061, id_1713, id_1716);
nand ( id_1071, id_1721, id_1724);
nand ( id_1103, id_1745, id_1748);
nand ( id_1115, id_1753, id_1756);
nand ( id_1157, id_1785, id_1788);
nand ( id_1169, id_1793, id_1796);
not ( id_1184, id_363);
nand ( id_1202, id_1197, id_1200);
nand ( id_1259, id_1841, id_1844);
nand ( id_1271, id_1849, id_1852);
not ( id_1322, id_406);
nand ( id_374, id_372, id_373);
nand ( id_396, id_1317, id_1320);
not ( id_1321, id_1317);
not ( id_1424, id_1418);
not ( id_1416, id_1410);
not ( id_1440, id_1434);
not ( id_1432, id_1426);
nand ( id_985, id_983, id_984);
nand ( id_995, id_993, id_994);
nand ( id_1035, id_1033, id_1034);
nand ( id_1045, id_1043, id_1044);
nand ( id_1063, id_1061, id_1062);
nand ( id_1073, id_1071, id_1072);
nand ( id_1105, id_1103, id_1104);
nand ( id_1117, id_1115, id_1116);
nand ( id_1159, id_1157, id_1158);
nand ( id_1171, id_1169, id_1170);
nand ( id_1212, id_1202, id_1203);
not ( id_1231, id_1227);
nand ( id_1232, id_1227, id_1230);
not ( id_1253, id_1249);
nand ( id_1254, id_1249, id_1252);
nand ( id_1261, id_1259, id_1260);
nand ( id_1273, id_1271, id_1272);
not ( id_1287, id_1283);
nand ( id_1288, id_1283, id_1286);
not ( id_1309, id_1305);
nand ( id_1310, id_1305, id_1308);
not ( id_1192, id_1184);
nand ( id_397, id_1312, id_1321);
not ( id_1330, id_1322);
buf ( id_1000, id_269);
buf ( id_1010, id_269);
nand ( id_1233, id_1222, id_1231);
nand ( id_1255, id_1244, id_1253);
nand ( id_1289, id_1278, id_1287);
nand ( id_1311, id_1300, id_1309);
not ( id_1381, id_374);
nand ( id_257, id_995, id_998);
not ( id_999, id_995);
nand ( id_260, id_985, id_988);
not ( id_989, id_985);
nand ( id_272, id_1035, id_1038);
not ( id_1039, id_1035);
nand ( id_294, id_1045, id_1048);
not ( id_1049, id_1045);
nand ( id_305, id_1073, id_1076);
not ( id_1077, id_1073);
nand ( id_308, id_1063, id_1066);
not ( id_1067, id_1063);
nand ( id_333, id_1117, id_1120);
not ( id_1121, id_1117);
nand ( id_358, id_1171, id_1174);
not ( id_1175, id_1171);
not ( id_1220, id_1212);
nand ( id_388, id_1273, id_1276);
not ( id_1277, id_1273);
nand ( id_398, id_396, id_397);
not ( id_1109, id_1105);
nand ( id_1110, id_1105, id_1108);
not ( id_1163, id_1159);
nand ( id_1164, id_1159, id_1162);
nand ( id_1234, id_1232, id_1233);
not ( id_1265, id_1261);
nand ( id_1266, id_1261, id_1264);
nand ( id_1822, id_1254, id_1255);
nand ( id_1862, id_1310, id_1311);
nand ( id_1865, id_1288, id_1289);
nand ( id_258, id_990, id_999);
nand ( id_261, id_980, id_989);
nand ( id_273, id_1030, id_1039);
not ( id_1018, id_1010);
not ( id_1008, id_1000);
nand ( id_295, id_1040, id_1049);
nand ( id_306, id_1068, id_1077);
nand ( id_309, id_1058, id_1067);
nand ( id_334, id_1112, id_1121);
nand ( id_359, id_1166, id_1175);
nand ( id_389, id_1268, id_1277);
not ( id_1385, id_1381);
nand ( id_1111, id_1100, id_1109);
nand ( id_1165, id_1154, id_1163);
nand ( id_1267, id_1256, id_1265);
not ( id_1886, id_398);
nand ( id_259, id_257, id_258);
nand ( id_262, id_260, id_261);
nand ( id_274, id_272, id_273);
nand ( id_296, id_294, id_295);
nand ( id_307, id_305, id_306);
nand ( id_310, id_308, id_309);
nand ( id_335, id_333, id_334);
nand ( id_360, id_358, id_359);
not ( id_1242, id_1234);
nand ( id_390, id_388, id_389);
not ( id_1828, id_1822);
not ( id_1868, id_1862);
not ( id_1869, id_1865);
nand ( id_1373, id_1164, id_1165);
nand ( id_1798, id_1110, id_1111);
nand ( id_1825, id_1266, id_1267);
not ( id_265, id_259);
not ( id_314, id_307);
not ( id_336, id_335);
not ( id_407, id_296);
nand ( id_1293, id_1865, id_1868);
nand ( id_1294, id_1862, id_1869);
not ( id_1892, id_1886);
not ( id_1777, id_360);
not ( id_1889, id_390);
buf ( id_410, id_310);
not ( id_1377, id_1373);
not ( id_1804, id_1798);
nand ( id_1237, id_1825, id_1828);
not ( id_1829, id_1825);
nand ( id_1295, id_1293, id_1294);
buf ( id_1670, id_274);
buf ( id_1678, id_274);
buf ( id_1729, id_310);
buf ( id_1737, id_310);
buf ( id_1761, id_262);
buf ( id_1769, id_262);
buf ( id_340, id_336);
buf ( id_343, id_314);
not ( id_1781, id_1777);
nand ( id_1238, id_1822, id_1829);
nand ( id_1325, id_1889, id_1892);
not ( id_1893, id_1889);
buf ( id_1340, id_407);
buf ( id_1352, id_407);
buf ( id_1673, id_265);
buf ( id_1681, id_265);
buf ( id_1801, id_314);
buf ( id_1897, id_336);
buf ( id_1905, id_336);
nand ( id_391, id_1295, id_1298);
not ( id_1299, id_1295);
not ( id_1676, id_1670);
not ( id_1684, id_1678);
nand ( id_1081, id_1729, id_1732);
not ( id_1733, id_1729);
nand ( id_1093, id_1737, id_1740);
not ( id_1741, id_1737);
not ( id_1765, id_1761);
not ( id_1773, id_1769);
nand ( id_1239, id_1237, id_1238);
nand ( id_1326, id_1886, id_1893);
buf ( id_1894, id_410);
buf ( id_1902, id_410);
nand ( id_392, id_1290, id_1299);
not ( id_1360, id_1352);
nand ( id_1003, id_1673, id_1676);
not ( id_1677, id_1673);
nand ( id_1013, id_1681, id_1684);
not ( id_1685, id_1681);
nand ( id_1082, id_1726, id_1733);
nand ( id_1094, id_1734, id_1741);
buf ( id_1122, id_340);
buf ( id_1134, id_340);
nand ( id_1187, id_1801, id_1804);
not ( id_1805, id_1801);
nand ( id_1327, id_1325, id_1326);
not ( id_1901, id_1897);
not ( id_1348, id_1340);
not ( id_1909, id_1905);
buf ( id_1758, id_343);
buf ( id_1766, id_343);
nand ( id_377, id_1239, id_1242);
not ( id_1243, id_1239);
nand ( id_393, id_391, id_392);
nand ( id_1004, id_1670, id_1677);
nand ( id_1014, id_1678, id_1685);
nand ( id_1083, id_1081, id_1082);
nand ( id_1095, id_1093, id_1094);
nand ( id_1188, id_1798, id_1805);
not ( id_1900, id_1894);
nand ( id_1344, id_1894, id_1901);
not ( id_1908, id_1902);
nand ( id_1356, id_1902, id_1909);
not ( id_1142, id_1134);
nand ( id_378, id_1234, id_1243);
nand ( id_399, id_1327, id_1330);
not ( id_1331, id_1327);
nand ( id_1005, id_1003, id_1004);
nand ( id_1015, id_1013, id_1014);
not ( id_1764, id_1758);
nand ( id_1126, id_1758, id_1765);
not ( id_1130, id_1122);
not ( id_1772, id_1766);
nand ( id_1138, id_1766, id_1773);
nand ( id_1189, id_1187, id_1188);
nand ( id_1343, id_1897, id_1900);
nand ( id_1355, id_1905, id_1908);
nand ( id_324, id_1095, id_1098);
not ( id_1099, id_1095);
nand ( id_379, id_377, id_378);
nand ( id_400, id_1322, id_1331);
nand ( id_449, id_393, id_918);
not ( id_1087, id_1083);
nand ( id_1088, id_1083, id_1086);
nand ( id_1125, id_1761, id_1764);
nand ( id_1137, id_1769, id_1772);
nand ( id_1345, id_1343, id_1344);
nand ( id_1357, id_1355, id_1356);
buf ( id_1397, id_393);
nand ( id_277, id_1015, id_1018);
not ( id_1019, id_1015);
nand ( id_280, id_1005, id_1008);
not ( id_1009, id_1005);
nand ( id_325, id_1090, id_1099);
nand ( id_364, id_1189, id_1192);
not ( id_1193, id_1189);
nand ( id_401, id_399, id_400);
nand ( id_1089, id_1078, id_1087);
nand ( id_1127, id_1125, id_1126);
nand ( id_1139, id_1137, id_1138);
nand ( id_278, id_1010, id_1019);
nand ( id_281, id_1000, id_1009);
nand ( id_326, id_324, id_325);
nand ( id_365, id_1184, id_1193);
nand ( id_413, id_1357, id_1360);
not ( id_1361, id_1357);
not ( id_1401, id_1397);
nand ( id_445, id_379, id_918);
not ( id_1349, id_1345);
nand ( id_1350, id_1345, id_1348);
buf ( id_1389, id_379);
buf ( id_1493, id_449);
buf ( id_1501, id_449);
nand ( id_1689, id_1088, id_1089);
nand ( id_279, id_277, id_278);
nand ( id_282, id_280, id_281);
nand ( id_346, id_1139, id_1142);
not ( id_1143, id_1139);
nand ( id_366, id_364, id_365);
nand ( id_414, id_1352, id_1361);
nand ( id_453, id_401, id_918);
not ( id_1131, id_1127);
nand ( id_1132, id_1127, id_1130);
nand ( id_1351, id_1340, id_1349);
not ( id_1365, id_326);
buf ( id_1405, id_401);
not ( id_285, id_279);
nand ( id_347, id_1134, id_1143);
not ( id_367, id_366);
nand ( id_415, id_413, id_414);
not ( id_1393, id_1389);
nand ( id_556, id_1501, id_1504);
not ( id_1505, id_1501);
nand ( id_559, id_1493, id_1496);
not ( id_1497, id_1493);
not ( id_1693, id_1689);
nand ( id_1133, id_1122, id_1131);
buf ( id_1477, id_445);
buf ( id_1485, id_445);
nand ( id_1809, id_1350, id_1351);
nand ( id_348, id_346, id_347);
not ( id_1369, id_1365);
not ( id_1409, id_1405);
nand ( id_557, id_1498, id_1505);
nand ( id_560, id_1490, id_1497);
buf ( id_1362, id_282);
not ( id_1378, id_415);
buf ( id_1429, id_453);
buf ( id_1437, id_453);
buf ( id_1686, id_282);
nand ( id_1774, id_1132, id_1133);
and ( id_1910, id_285, id_853);
and ( id_1918, id_856, id_367);
nand ( id_544, id_1485, id_1488);
not ( id_1489, id_1485);
nand ( id_547, id_1477, id_1480);
not ( id_1481, id_1477);
nand ( id_558, id_556, id_557);
nand ( id_561, id_559, id_560);
not ( id_1813, id_1809);
not ( id_1370, id_348);
not ( id_1368, id_1362);
nand ( id_417, id_1362, id_1369);
not ( id_1384, id_1378);
nand ( id_424, id_1378, id_1385);
nand ( id_508, id_1437, id_1440);
not ( id_1441, id_1437);
nand ( id_511, id_1429, id_1432);
not ( id_1433, id_1429);
nand ( id_545, id_1482, id_1489);
nand ( id_548, id_1474, id_1481);
not ( id_564, id_558);
not ( id_1692, id_1686);
nand ( id_1024, id_1686, id_1693);
not ( id_1780, id_1774);
nand ( id_1148, id_1774, id_1781);
not ( id_1916, id_1910);
not ( id_1924, id_1918);
nand ( id_416, id_1365, id_1368);
not ( id_1376, id_1370);
nand ( id_421, id_1370, id_1377);
nand ( id_423, id_1381, id_1384);
nand ( id_509, id_1434, id_1441);
nand ( id_512, id_1426, id_1433);
nand ( id_546, id_544, id_545);
nand ( id_549, id_547, id_548);
not ( id_719, id_561);
buf ( id_722, id_561);
nand ( id_1023, id_1689, id_1692);
nand ( id_1147, id_1777, id_1780);
nand ( id_418, id_416, id_417);
nand ( id_420, id_1373, id_1376);
nand ( id_425, id_423, id_424);
nand ( id_510, id_508, id_509);
nand ( id_513, id_511, id_512);
not ( id_552, id_546);
nand ( id_1025, id_1023, id_1024);
nand ( id_1149, id_1147, id_1148);
not ( id_419, id_418);
nand ( id_422, id_420, id_421);
nand ( id_441, id_425, id_918);
not ( id_516, id_510);
not ( id_725, id_549);
buf ( id_728, id_549);
not ( id_1029, id_1025);
not ( id_1153, id_1149);
nand ( id_433, id_419, id_918);
nand ( id_437, id_422, id_918);
not ( id_663, id_513);
buf ( id_666, id_513);
and ( id_731, id_719, id_725);
and ( id_746, id_722, id_725);
and ( id_756, id_719, id_728);
and ( id_770, id_722, id_728);
buf ( id_1461, id_441);
buf ( id_1469, id_441);
buf ( id_1413, id_433);
buf ( id_1421, id_433);
buf ( id_1445, id_437);
buf ( id_1453, id_437);
nand ( id_532, id_1469, id_1472);
not ( id_1473, id_1469);
nand ( id_535, id_1461, id_1464);
not ( id_1465, id_1461);
nand ( id_495, id_1421, id_1424);
not ( id_1425, id_1421);
nand ( id_498, id_1413, id_1416);
not ( id_1417, id_1413);
nand ( id_520, id_1453, id_1456);
not ( id_1457, id_1453);
nand ( id_523, id_1445, id_1448);
not ( id_1449, id_1445);
nand ( id_533, id_1466, id_1473);
nand ( id_536, id_1458, id_1465);
nand ( id_496, id_1418, id_1425);
nand ( id_499, id_1410, id_1417);
nand ( id_521, id_1450, id_1457);
nand ( id_524, id_1442, id_1449);
nand ( id_534, id_532, id_533);
nand ( id_537, id_535, id_536);
nand ( id_497, id_495, id_496);
nand ( id_500, id_498, id_499);
nand ( id_522, id_520, id_521);
nand ( id_525, id_523, id_524);
not ( id_540, id_534);
not ( id_503, id_497);
not ( id_528, id_522);
not ( id_669, id_537);
buf ( id_672, id_537);
not ( id_569, id_500);
and ( id_588, id_566, id_500);
not ( id_618, id_525);
and ( id_639, id_615, id_525);
nand ( id_867, id_516, id_564, id_552, id_540, id_482, id_528, id_503, id_487);
buf ( id_588a, id_588);
buf ( id_588b, id_588);
buf ( id_639a, id_639);
buf ( id_639b, id_639);
and ( id_675, id_663, id_669);
and ( id_688, id_666, id_669);
and ( id_696, id_663, id_672);
and ( id_710, id_666, id_672);
and ( id_73, id_949, id_867, id_932);
buf ( id_572, id_569);
and ( id_573, id_566, id_569);
buf ( id_621, id_618);
and ( id_622, id_615, id_618);
nand ( id_776, id_588a, id_639a, id_696, id_731, id_958);
nand ( id_780, id_588a, id_639a, id_675, id_756, id_958);
nand ( id_784, id_588a, id_639a, id_675, id_746, id_958);
nand ( id_788, id_588a, id_639a, id_688, id_731, id_958);
nand ( id_812, id_588b, id_639a, id_710, id_746, id_969);
nand ( id_832, id_588b, id_639b, id_696, id_770, id_969);
nand ( id_836, id_588b, id_639b, id_710, id_756, id_969);
and ( id_1509, id_588a, id_639a, id_696, id_731, id_958);
and ( id_1517, id_588a, id_639a, id_675, id_756, id_958);
and ( id_1525, id_588a, id_639a, id_675, id_746, id_958);
and ( id_1533, id_588a, id_639a, id_688, id_731, id_958);
and ( id_1581, id_588b, id_639a, id_710, id_746, id_969);
and ( id_1621, id_588b, id_639b, id_696, id_770, id_969);
and ( id_1629, id_588b, id_639b, id_710, id_756, id_969);
nand ( id_792, id_588a, id_622, id_696, id_756, id_958);
nand ( id_796, id_588b, id_622, id_696, id_746, id_958);
nand ( id_800, id_588b, id_622, id_710, id_731, id_958);
nand ( id_804, id_588b, id_622, id_675, id_770, id_958);
nand ( id_808, id_588b, id_622, id_688, id_756, id_969);
nand ( id_816, id_573, id_639b, id_696, id_756, id_969);
nand ( id_820, id_573, id_639b, id_696, id_746, id_969);
nand ( id_824, id_573, id_639b, id_710, id_731, id_969);
nand ( id_828, id_573, id_639b, id_688, id_756, id_969);
nand ( id_871, id_588b, id_622, id_675, id_731, id_979);
nand ( id_873, id_573, id_639b, id_675, id_731, id_979);
nand ( id_875, id_573, id_622, id_696, id_731, id_979);
nand ( id_877, id_573, id_622, id_675, id_756, id_979);
nand ( id_879, id_573, id_622, id_675, id_746, id_979);
nand ( id_881, id_573, id_622, id_688, id_731, id_979);
nand ( id_883, id_573, id_621, id_675, id_731, id_979);
nand ( id_885, id_572, id_622, id_675, id_731, id_979);
and ( id_1541, id_588a, id_622, id_696, id_756, id_958);
and ( id_1549, id_588b, id_622, id_696, id_746, id_958);
and ( id_1557, id_588b, id_622, id_710, id_731, id_958);
and ( id_1565, id_588b, id_622, id_675, id_770, id_958);
and ( id_1573, id_588b, id_622, id_688, id_756, id_969);
and ( id_1589, id_573, id_639b, id_696, id_756, id_969);
and ( id_1597, id_573, id_639b, id_696, id_746, id_969);
and ( id_1605, id_573, id_639b, id_710, id_731, id_969);
and ( id_1613, id_573, id_639b, id_688, id_756, id_969);
nand ( id_1, id_1509, id_1512);
not ( id_1513, id_1509);
nand ( id_4, id_1517, id_1520);
not ( id_1521, id_1517);
nand ( id_7, id_1525, id_1528);
not ( id_1529, id_1525);
nand ( id_10, id_1533, id_1536);
not ( id_1537, id_1533);
nand ( id_28, id_1581, id_1584);
not ( id_1585, id_1581);
nand ( id_43, id_1621, id_1624);
not ( id_1625, id_1621);
nand ( id_46, id_1629, id_1632);
not ( id_1633, id_1629);
and ( id_886, id_871, id_873, id_875, id_877, id_879, id_881, id_883, id_885);
nand ( id_2, id_1506, id_1513);
nand ( id_5, id_1514, id_1521);
nand ( id_8, id_1522, id_1529);
nand ( id_11, id_1530, id_1537);
nand ( id_13, id_1541, id_1544);
not ( id_1545, id_1541);
nand ( id_16, id_1549, id_1552);
not ( id_1553, id_1549);
nand ( id_19, id_1557, id_1560);
not ( id_1561, id_1557);
nand ( id_22, id_1565, id_1568);
not ( id_1569, id_1565);
nand ( id_25, id_1573, id_1576);
not ( id_1577, id_1573);
nand ( id_29, id_1578, id_1585);
nand ( id_31, id_1589, id_1592);
not ( id_1593, id_1589);
nand ( id_34, id_1597, id_1600);
not ( id_1601, id_1597);
nand ( id_37, id_1605, id_1608);
not ( id_1609, id_1605);
nand ( id_40, id_1613, id_1616);
not ( id_1617, id_1613);
nand ( id_44, id_1618, id_1625);
nand ( id_47, id_1626, id_1633);
nand ( id_857, id_776, id_780, id_784, id_788, id_792, id_796, id_800, id_804);
nand ( id_860, id_808, id_812, id_816, id_820, id_824, id_828, id_832, id_836);
and ( id_863, id_776, id_780, id_784, id_788, id_792, id_796, id_800, id_804);
and ( id_865, id_808, id_812, id_816, id_820, id_824, id_828, id_832, id_836);
nand ( id_3, id_1, id_2);
nand ( id_6, id_4, id_5);
nand ( id_9, id_7, id_8);
nand ( id_12, id_10, id_11);
nand ( id_14, id_1538, id_1545);
nand ( id_17, id_1546, id_1553);
nand ( id_20, id_1554, id_1561);
nand ( id_23, id_1562, id_1569);
nand ( id_26, id_1570, id_1577);
nand ( id_30, id_28, id_29);
nand ( id_32, id_1586, id_1593);
nand ( id_35, id_1594, id_1601);
nand ( id_38, id_1602, id_1609);
nand ( id_41, id_1610, id_1617);
nand ( id_45, id_43, id_44);
nand ( id_48, id_46, id_47);
and ( id_1913, id_857, id_859);
and ( id_1921, id_860, id_862);
nand ( id_15, id_13, id_14);
nand ( id_18, id_16, id_17);
nand ( id_21, id_19, id_20);
nand ( id_24, id_22, id_23);
nand ( id_27, id_25, id_26);
nand ( id_33, id_31, id_32);
nand ( id_36, id_34, id_35);
nand ( id_39, id_37, id_38);
nand ( id_42, id_40, id_41);
and ( id_887, id_863, id_865, id_886);
nand ( id_462, id_863, id_865);
and ( id_74, id_949, id_867, id_887);
nand ( id_1637, id_1913, id_1916);
not ( id_1917, id_1913);
nand ( id_1647, id_1921, id_1924);
not ( id_1925, id_1921);
nor ( id_75, id_73, id_74);
and ( id_1020, id_457, id_911, id_462);
and ( id_1144, id_469, id_911, id_462);
and ( id_1386, id_475, id_911, id_462);
and ( id_1394, id_478, id_911, id_462);
and ( id_1402, id_459, id_911, id_462);
nand ( id_1638, id_1910, id_1917);
nand ( id_1648, id_1918, id_1925);
and ( id_1806, id_472, id_911, id_462);
nand ( id_1639, id_1637, id_1638);
nand ( id_1649, id_1647, id_1648);
nand ( id_287, id_1020, id_1029);
nand ( id_350, id_1144, id_1153);
nand ( id_427, id_1386, id_1393);
nand ( id_429, id_1394, id_1401);
nand ( id_431, id_1402, id_1409);
not ( id_1028, id_1020);
not ( id_1152, id_1144);
not ( id_1392, id_1386);
not ( id_1400, id_1394);
not ( id_1408, id_1402);
not ( id_1812, id_1806);
nand ( id_1216, id_1806, id_1813);
nand ( id_286, id_1025, id_1028);
nand ( id_349, id_1149, id_1152);
nand ( id_426, id_1389, id_1392);
nand ( id_428, id_1397, id_1400);
nand ( id_430, id_1405, id_1408);
nand ( id_67, id_1639, id_1642);
not ( id_1643, id_1639);
nand ( id_70, id_1649, id_1652);
not ( id_1653, id_1649);
nand ( id_1215, id_1809, id_1812);
nand ( id_49, id_286, id_287);
nand ( id_53, id_349, id_350);
nand ( id_59, id_426, id_427);
nand ( id_61, id_428, id_429);
nand ( id_65, id_430, id_431);
nand ( id_68, id_1634, id_1643);
nand ( id_71, id_1644, id_1653);
nand ( id_1217, id_1215, id_1216);
and ( id_51, id_49, id_50);
and ( id_54, id_52, id_53);
and ( id_60, id_58, id_59);
and ( id_63, id_61, id_62);
and ( id_66, id_64, id_65);
nand ( id_69, id_67, id_68);
nand ( id_72, id_70, id_71);
nand ( id_375, id_1217, id_1220);
not ( id_1221, id_1217);
nand ( id_376, id_1212, id_1221);
nand ( id_55, id_375, id_376);
and ( id_57, id_55, id_56);

endmodule
