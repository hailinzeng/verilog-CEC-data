module c3540
( id_1 ,id_13 ,id_20 ,id_33 ,id_41 ,id_45 ,id_50 ,id_58 ,id_68 ,id_77 ,id_87 ,id_97 ,id_107 ,id_116 ,id_124 ,id_125 ,id_128 ,id_132 ,id_137 ,id_143 ,id_150 ,id_159 ,id_169 ,id_179 ,id_190 ,id_200 ,id_213 ,id_222 ,id_223 ,id_226 ,id_232 ,id_238 ,id_244 ,id_250 ,id_257 ,id_264 ,id_270 ,id_274 ,id_283 ,id_294 ,id_303 ,id_311 ,id_317 ,id_322 ,id_326 ,id_329 ,id_330 ,id_343 ,id_1698 ,id_2897 ,id_353 ,id_355 ,id_361 ,id_358 ,id_351 ,id_372 ,id_369 ,id_399 ,id_364 ,id_396 ,id_384 ,id_367 ,id_387 ,id_393 ,id_390 ,id_378 ,id_375 ,id_381 ,id_407 ,id_409 ,id_405 ,id_402 );

input id_1, id_13, id_20, id_33, id_41, id_45, id_50, id_58, id_68, id_77, id_87, id_97, id_107, id_116, id_124, id_125, id_128, id_132, id_137, id_143, id_150, id_159, id_169, id_179, id_190, id_200, id_213, id_222, id_223, id_226, id_232, id_238, id_244, id_250, id_257, id_264, id_270, id_274, id_283, id_294, id_303, id_311, id_317, id_322, id_326, id_329, id_330, id_343, id_1698, id_2897;

output id_353, id_355, id_361, id_358, id_351, id_372, id_369, id_399, id_364, id_396, id_384, id_367, id_387, id_393, id_390, id_378, id_375, id_381, id_407, id_409, id_405, id_402;

buf ( id_432, id_50);
not ( id_442, id_50);
buf ( id_447, id_58);
not ( id_456, id_58);
buf ( id_460, id_68);
not ( id_463, id_68);
buf ( id_467, id_68);
buf ( id_476, id_77);
not ( id_479, id_77);
buf ( id_483, id_77);
buf ( id_492, id_87);
not ( id_501, id_87);
buf ( id_504, id_97);
not ( id_513, id_97);
buf ( id_517, id_107);
not ( id_526, id_107);
buf ( id_530, id_116);
not ( id_540, id_116);
or ( id_587, id_257, id_264);
not ( id_704, id_1);
buf ( id_707, id_1);
not ( id_714, id_1);
buf ( id_717, id_13);
not ( id_724, id_13);
and ( id_731, id_13, id_20);
not ( id_732, id_20);
buf ( id_736, id_20);
not ( id_741, id_20);
not ( id_758, id_33);
buf ( id_776, id_33);
not ( id_780, id_33);
and ( id_788, id_33, id_41);
not ( id_791, id_41);
or ( id_798, id_41, id_45);
buf ( id_799, id_45);
not ( id_802, id_45);
not ( id_826, id_50);
buf ( id_828, id_58);
not ( id_831, id_58);
buf ( id_833, id_68);
not ( id_836, id_68);
buf ( id_839, id_87);
not ( id_842, id_87);
buf ( id_845, id_97);
not ( id_848, id_97);
not ( id_851, id_107);
buf ( id_890, id_1);
buf ( id_898, id_68);
buf ( id_907, id_107);
not ( id_1032, id_20);
buf ( id_1035, id_190);
not ( id_1048, id_200);
and ( id_1049, id_20, id_200);
nand ( id_1050, id_20, id_200);
and ( id_1051, id_20, id_179);
not ( id_1540, id_20);
or ( id_1699, id_1698, id_33);
nand ( id_1826, id_1, id_13);
nand ( id_1827, id_1, id_20, id_33);
not ( id_1828, id_20);
not ( id_2051, id_33);
buf ( id_2478, id_179);
not ( id_2865, id_213);
buf ( id_2868, id_343);
buf ( id_2931, id_226);
buf ( id_2934, id_232);
buf ( id_2939, id_238);
buf ( id_2942, id_244);
buf ( id_2947, id_250);
buf ( id_2950, id_257);
buf ( id_2957, id_264);
buf ( id_2960, id_270);
buf ( id_3007, id_50);
buf ( id_3079, id_58);
buf ( id_3087, id_58);
buf ( id_3095, id_97);
buf ( id_3103, id_97);
buf ( id_3419, id_330);
and ( id_588, id_250, id_587);
or ( id_759, id_758, id_20);
or ( id_1541, id_1540, id_169);
not ( id_1772, id_731);
or ( id_1829, id_1828, id_1);
and ( id_1834, id_1826, id_1827);
or ( id_2052, id_2051, id_1);
and ( id_625, id_826, id_831, id_836);
nand ( id_545, id_226, id_432);
nand ( id_546, id_232, id_447);
nand ( id_547, id_238, id_467);
nand ( id_548, id_244, id_483);
nand ( id_549, id_250, id_492);
nand ( id_550, id_257, id_504);
nand ( id_551, id_264, id_517);
nand ( id_552, id_270, id_530);
not ( id_2937, id_2931);
not ( id_2938, id_2934);
not ( id_2945, id_2939);
not ( id_2946, id_2942);
nand ( id_621, id_456, id_463);
nand ( id_626, id_513, id_526);
nand ( id_635, id_460, id_476);
buf ( id_636, id_442);
not ( id_3085, id_3079);
not ( id_3101, id_3095);
buf ( id_657, id_802);
buf ( id_675, id_802);
buf ( id_721, id_717);
buf ( id_784, id_780);
buf ( id_794, id_791);
and ( id_807, id_714, id_798);
and ( id_816, id_714, id_799, id_791);
and ( id_823, id_704, id_799);
and ( id_860, id_707, id_724, id_736);
nand ( id_861, id_707, id_724, id_736);
nand ( id_864, id_707, id_724);
buf ( id_893, id_890);
nand ( id_896, id_717, id_732, id_45);
nand ( id_897, id_826, id_831, id_836);
not ( id_3093, id_3087);
and ( id_905, id_842, id_848, id_851);
nand ( id_906, id_842, id_848, id_851);
not ( id_3109, id_3103);
not ( id_973, id_741);
not ( id_980, id_741);
not ( id_987, id_741);
not ( id_994, id_741);
not ( id_1001, id_741);
not ( id_1008, id_741);
not ( id_1015, id_741);
not ( id_1022, id_741);
or ( id_1038, id_1032, id_1035);
nor ( id_1043, id_1032, id_1035);
buf ( id_1054, id_1051);
not ( id_1057, id_1051);
buf ( id_1512, id_776);
buf ( id_1681, id_780);
not ( id_1717, id_1699);
not ( id_1724, id_1699);
not ( id_1731, id_1699);
not ( id_1738, id_1699);
not ( id_1745, id_1699);
not ( id_1752, id_1699);
not ( id_1759, id_1699);
not ( id_1766, id_1699);
or ( id_1773, id_1, id_1772);
not ( id_1790, id_788);
not ( id_1808, id_788);
and ( id_2278, id_704, id_717, id_732);
not ( id_2481, id_2478);
not ( id_3425, id_3419);
or ( id_2871, id_2865, id_2868);
nor ( id_2874, id_2865, id_2868);
not ( id_2953, id_2947);
not ( id_2954, id_2950);
not ( id_2963, id_2957);
not ( id_2964, id_2960);
buf ( id_3010, id_456);
not ( id_3013, id_3007);
buf ( id_3017, id_463);
buf ( id_3020, id_479);
buf ( id_3027, id_501);
buf ( id_3030, id_513);
buf ( id_3037, id_526);
buf ( id_3040, id_540);
buf ( id_3082, id_898);
buf ( id_3090, id_898);
buf ( id_3098, id_907);
buf ( id_3106, id_907);
nand ( id_352, id_479, id_625);
and ( id_553, id_545, id_546, id_547, id_548);
and ( id_554, id_549, id_550, id_551, id_552);
nand ( id_555, id_2934, id_2937);
nand ( id_556, id_2931, id_2938);
nand ( id_560, id_2942, id_2945);
nand ( id_561, id_2939, id_2946);
and ( id_650, id_432, id_621);
and ( id_956, id_890, id_896);
not ( id_974, id_759);
and ( id_975, id_741, id_759);
and ( id_976, id_897, id_973);
not ( id_981, id_759);
and ( id_982, id_741, id_759);
not ( id_988, id_759);
and ( id_989, id_741, id_759);
and ( id_990, id_836, id_987);
not ( id_995, id_759);
and ( id_996, id_741, id_759);
and ( id_997, id_77, id_994);
not ( id_1002, id_759);
and ( id_1003, id_741, id_759);
and ( id_1004, id_906, id_1001);
not ( id_1009, id_759);
and ( id_1010, id_741, id_759);
not ( id_1016, id_759);
and ( id_1017, id_741, id_759);
and ( id_1018, id_851, id_1015);
not ( id_1023, id_759);
and ( id_1024, id_741, id_759);
and ( id_1025, id_116, id_1022);
and ( id_1720, id_222, id_1717);
and ( id_1727, id_223, id_1724);
and ( id_1734, id_226, id_1731);
and ( id_1741, id_232, id_1738);
and ( id_1748, id_238, id_1745);
and ( id_1755, id_244, id_1752);
and ( id_1762, id_250, id_1759);
and ( id_1769, id_257, id_1766);
and ( id_1791, id_1, id_13, id_1790);
and ( id_1809, id_1, id_13, id_1808);
not ( id_1851, id_1834);
not ( id_1901, id_1834);
not ( id_1952, id_1834);
not ( id_2002, id_1834);
not ( id_2057, id_1834);
not ( id_2109, id_1834);
not ( id_2162, id_1834);
not ( id_2214, id_1834);
nand ( id_2955, id_2950, id_2953);
nand ( id_2956, id_2947, id_2954);
nand ( id_2965, id_2960, id_2963);
nand ( id_2966, id_2957, id_2964);
not ( id_353, id_352);
and ( id_354, id_87, id_626);
nand ( id_557, id_555, id_556);
nand ( id_562, id_560, id_561);
nand ( id_586, id_553, id_554);
and ( id_630, id_540, id_905);
nand ( id_634, id_540, id_905);
not ( id_639, id_636);
nand ( id_642, id_3082, id_3085);
not ( id_3086, id_3082);
and ( id_644, id_460, id_636);
nand ( id_646, id_3098, id_3101);
not ( id_3102, id_3098);
nand ( id_654, id_87, id_626);
not ( id_660, id_657);
not ( id_678, id_675);
nand ( id_804, id_860, id_776);
nand ( id_806, id_860, id_780);
nand ( id_855, id_707, id_721, id_736);
nand ( id_867, id_707, id_724, id_736, id_794);
nand ( id_903, id_3090, id_3093);
not ( id_3094, id_3090);
nand ( id_912, id_3106, id_3109);
not ( id_3110, id_3106);
not ( id_915, id_861);
not ( id_927, id_893);
not ( id_941, id_864);
and ( id_977, id_828, id_974);
and ( id_978, id_150, id_975);
and ( id_984, id_833, id_981);
and ( id_985, id_159, id_982);
and ( id_991, id_77, id_988);
and ( id_992, id_50, id_989);
and ( id_998, id_839, id_995);
and ( id_999, id_828, id_996);
and ( id_1005, id_845, id_1002);
and ( id_1006, id_833, id_1003);
and ( id_1012, id_107, id_1009);
and ( id_1013, id_77, id_1010);
and ( id_1019, id_116, id_1016);
and ( id_1020, id_839, id_1017);
and ( id_1026, id_283, id_1023);
and ( id_1027, id_845, id_1024);
and ( id_1060, id_200, id_1054);
and ( id_1063, id_1048, id_1054);
and ( id_1066, id_1049, id_1057);
and ( id_1069, id_1050, id_1057);
nand ( id_1527, id_784, id_794);
nand ( id_1530, id_776, id_794);
nand ( id_1542, id_707, id_721, id_1541);
nand ( id_1563, id_724, id_732, id_784);
nand ( id_1572, id_724, id_784);
not ( id_1581, id_1512);
not ( id_1585, id_1512);
not ( id_1589, id_1512);
not ( id_1593, id_1512);
not ( id_1597, id_1512);
not ( id_1601, id_1512);
not ( id_1605, id_1512);
not ( id_1716, id_1681);
and ( id_1718, id_1681, id_1699);
not ( id_1723, id_1681);
and ( id_1725, id_1681, id_1699);
not ( id_1730, id_1681);
and ( id_1732, id_1681, id_1699);
not ( id_1737, id_1681);
and ( id_1739, id_1681, id_1699);
not ( id_1744, id_1681);
and ( id_1746, id_1681, id_1699);
not ( id_1751, id_1681);
and ( id_1753, id_1681, id_1699);
not ( id_1758, id_1681);
and ( id_1760, id_1681, id_1699);
not ( id_1765, id_1681);
and ( id_1767, id_1681, id_1699);
and ( id_1852, id_1834, id_1773);
nor ( id_1856, id_50, id_1773);
not ( id_1870, id_807);
and ( id_1902, id_1834, id_1773);
nor ( id_1906, id_58, id_1773);
not ( id_1920, id_807);
and ( id_1953, id_1834, id_1773);
nor ( id_1957, id_68, id_1773);
not ( id_1971, id_807);
and ( id_2003, id_1834, id_1773);
nor ( id_2007, id_77, id_1773);
not ( id_2021, id_807);
and ( id_2058, id_1834, id_1773);
nor ( id_2062, id_87, id_1773);
not ( id_2076, id_823);
and ( id_2110, id_1834, id_1773);
nor ( id_2114, id_97, id_1773);
not ( id_2128, id_816);
and ( id_2163, id_1834, id_1773);
nor ( id_2167, id_107, id_1773);
not ( id_2181, id_816);
and ( id_2215, id_1834, id_1773);
nor ( id_2219, id_116, id_1773);
not ( id_2233, id_816);
and ( id_2285, id_2278, id_213);
nand ( id_2288, id_2278, id_213);
and ( id_2289, id_2278, id_213, id_343);
nand ( id_2293, id_2278, id_213, id_343);
and ( id_2298, id_2278, id_213, id_343);
nand ( id_2302, id_2278, id_213, id_343);
buf ( id_2877, id_2874);
nand ( id_2983, id_2955, id_2956);
nand ( id_2986, id_2965, id_2966);
not ( id_3014, id_3010);
nand ( id_3015, id_3010, id_3013);
not ( id_3023, id_3017);
not ( id_3024, id_3020);
not ( id_3033, id_3027);
not ( id_3034, id_3030);
not ( id_3043, id_3037);
not ( id_3044, id_3040);
not ( id_355, id_354);
nand ( id_643, id_3079, id_3086);
nand ( id_647, id_3095, id_3102);
and ( id_680, id_650, id_675);
nand ( id_904, id_3087, id_3094);
nand ( id_913, id_3103, id_3110);
and ( id_920, id_588, id_915);
or ( id_979, id_976, id_977, id_978);
or ( id_993, id_990, id_991, id_992);
or ( id_1000, id_997, id_998, id_999);
or ( id_1007, id_1004, id_1005, id_1006);
or ( id_1021, id_1018, id_1019, id_1020);
or ( id_1028, id_1025, id_1026, id_1027);
and ( id_1719, id_77, id_1716);
and ( id_1721, id_223, id_1718);
and ( id_1726, id_87, id_1723);
and ( id_1728, id_226, id_1725);
and ( id_1733, id_97, id_1730);
and ( id_1735, id_232, id_1732);
and ( id_1740, id_107, id_1737);
and ( id_1742, id_238, id_1739);
and ( id_1747, id_116, id_1744);
and ( id_1749, id_244, id_1746);
and ( id_1754, id_283, id_1751);
and ( id_1756, id_250, id_1753);
and ( id_1761, id_294, id_1758);
and ( id_1763, id_257, id_1760);
and ( id_1768, id_303, id_1765);
and ( id_1770, id_264, id_1767);
buf ( id_1794, id_1791);
not ( id_1799, id_1791);
buf ( id_1812, id_1809);
not ( id_1817, id_1809);
and ( id_1859, id_50, id_1829, id_1852);
and ( id_1909, id_58, id_1829, id_1902);
and ( id_1960, id_68, id_1829, id_1953);
and ( id_2010, id_77, id_1829, id_2003);
and ( id_2065, id_87, id_2052, id_2058);
and ( id_2117, id_97, id_2052, id_2110);
and ( id_2170, id_107, id_2052, id_2163);
and ( id_2222, id_116, id_2052, id_2215);
not ( id_2678, id_956);
not ( id_2697, id_956);
not ( id_2716, id_956);
not ( id_2733, id_956);
not ( id_2751, id_956);
not ( id_2768, id_956);
not ( id_2785, id_956);
not ( id_2802, id_956);
nand ( id_3016, id_3007, id_3014);
nand ( id_3025, id_3020, id_3023);
nand ( id_3026, id_3017, id_3024);
nand ( id_3035, id_3030, id_3033);
nand ( id_3036, id_3027, id_3034);
nand ( id_3045, id_3040, id_3043);
nand ( id_3046, id_3037, id_3044);
not ( id_2989, id_2983);
not ( id_2990, id_2986);
not ( id_610, id_804);
and ( id_613, id_804, id_806);
not ( id_616, id_806);
nand ( id_640, id_642, id_643);
nand ( id_648, id_646, id_647);
and ( id_655, id_630, id_635, id_442, id_58);
not ( id_665, id_804);
and ( id_668, id_804, id_806);
not ( id_671, id_806);
not ( id_683, id_804);
not ( id_685, id_806);
and ( id_688, id_804, id_806);
not ( id_694, id_804);
not ( id_696, id_806);
and ( id_699, id_804, id_806);
buf ( id_870, id_867);
buf ( id_887, id_867);
nand ( id_901, id_903, id_904);
nand ( id_910, id_912, id_913);
not ( id_914, id_855);
and ( id_916, id_855, id_861);
not ( id_942, id_855);
and ( id_943, id_864, id_855);
nand ( id_1072, id_1043, id_1069);
nand ( id_1084, id_1043, id_1066);
nand ( id_1096, id_1038, id_1069);
nand ( id_1108, id_1038, id_1066);
nand ( id_1120, id_1043, id_1063);
nand ( id_1132, id_1043, id_1060);
nand ( id_1144, id_1038, id_1063);
nand ( id_1156, id_1038, id_1060);
not ( id_1533, id_1527);
not ( id_1534, id_1530);
and ( id_1535, id_1527, id_1530);
buf ( id_1545, id_1542);
buf ( id_1554, id_1542);
not ( id_1610, id_1572);
not ( id_1619, id_1572);
not ( id_1628, id_1572);
not ( id_1637, id_1572);
not ( id_1646, id_1563);
not ( id_1655, id_1563);
not ( id_1664, id_1563);
not ( id_1673, id_1563);
or ( id_1722, id_1719, id_1720, id_1721);
or ( id_1729, id_1726, id_1727, id_1728);
or ( id_1736, id_1733, id_1734, id_1735);
or ( id_1743, id_1740, id_1741, id_1742);
or ( id_1750, id_1747, id_1748, id_1749);
or ( id_1757, id_1754, id_1755, id_1756);
or ( id_1764, id_1761, id_1762, id_1763);
or ( id_1771, id_1768, id_1769, id_1770);
and ( id_1853, id_979, id_1851);
and ( id_1954, id_993, id_1952);
and ( id_2004, id_1000, id_2002);
and ( id_2059, id_1007, id_2057);
and ( id_2164, id_1021, id_2162);
and ( id_2216, id_1028, id_2214);
buf ( id_2485, id_2293);
and ( id_2900, id_2877, id_2897);
nand ( id_2903, id_2877, id_2897);
buf ( id_2967, id_557);
buf ( id_2970, id_562);
buf ( id_2975, id_557);
buf ( id_2978, id_562);
nand ( id_3047, id_3015, id_3016);
nand ( id_3050, id_3025, id_3026);
nand ( id_3055, id_3035, id_3036);
nand ( id_3058, id_3045, id_3046);
nand ( id_574, id_2986, id_2989);
nand ( id_575, id_2983, id_2990);
and ( id_617, id_501, id_613);
and ( id_641, id_640, id_476, id_639);
and ( id_649, id_530, id_648);
and ( id_662, id_655, id_657);
and ( id_672, id_513, id_668);
and ( id_690, id_654, id_685);
and ( id_691, id_540, id_688);
and ( id_701, id_634, id_696);
and ( id_702, id_526, id_699);
not ( id_902, id_901);
not ( id_911, id_910);
and ( id_917, id_650, id_914);
and ( id_923, id_586, id_916);
and ( id_1538, id_442, id_1535);
and ( id_1871, id_1817, id_226, id_1870);
and ( id_1872, id_1817, id_274, id_807);
and ( id_1873, id_1812, id_1722);
and ( id_1921, id_1817, id_232, id_1920);
and ( id_1922, id_1817, id_274, id_807);
and ( id_1923, id_1812, id_1729);
and ( id_1972, id_1817, id_238, id_1971);
and ( id_1973, id_1817, id_274, id_807);
and ( id_1974, id_1812, id_1736);
and ( id_2022, id_1817, id_244, id_2021);
and ( id_2023, id_1817, id_274, id_807);
and ( id_2024, id_1812, id_1743);
and ( id_2077, id_1799, id_250, id_2076);
and ( id_2078, id_1799, id_274, id_823);
and ( id_2079, id_1794, id_1750);
and ( id_2129, id_1799, id_257, id_2128);
and ( id_2130, id_1799, id_274, id_816);
and ( id_2131, id_1794, id_1757);
and ( id_2182, id_1799, id_264, id_2181);
and ( id_2183, id_1799, id_274, id_816);
and ( id_2184, id_1794, id_1764);
and ( id_2234, id_1799, id_270, id_2233);
and ( id_2235, id_1799, id_274, id_816);
and ( id_2236, id_1794, id_1771);
not ( id_2973, id_2967);
not ( id_2974, id_2970);
not ( id_2981, id_2975);
not ( id_2982, id_2978);
nand ( id_576, id_574, id_575);
not ( id_3053, id_3047);
not ( id_3054, id_3050);
not ( id_3061, id_3055);
not ( id_3062, id_3058);
or ( id_645, id_641, id_644);
not ( id_926, id_887);
and ( id_928, id_887, id_893);
and ( id_947, id_649, id_942);
and ( id_983, id_902, id_980);
and ( id_1011, id_911, id_1008);
buf ( id_1075, id_1072);
buf ( id_1087, id_1084);
buf ( id_1099, id_1096);
buf ( id_1111, id_1108);
buf ( id_1123, id_1120);
buf ( id_1135, id_1132);
buf ( id_1147, id_1144);
buf ( id_1159, id_1156);
buf ( id_1168, id_1072);
buf ( id_1177, id_1084);
buf ( id_1186, id_1096);
buf ( id_1195, id_1108);
buf ( id_1204, id_1120);
buf ( id_1213, id_1132);
buf ( id_1222, id_1144);
buf ( id_1231, id_1156);
not ( id_1609, id_1545);
and ( id_1611, id_1545, id_1572);
not ( id_1618, id_1545);
and ( id_1620, id_1545, id_1572);
not ( id_1627, id_1545);
and ( id_1629, id_1545, id_1572);
not ( id_1636, id_1545);
and ( id_1638, id_1545, id_1572);
not ( id_1645, id_1554);
and ( id_1647, id_1554, id_1563);
not ( id_1654, id_1554);
and ( id_1656, id_1554, id_1563);
not ( id_1663, id_1554);
and ( id_1665, id_1554, id_1563);
not ( id_1672, id_1554);
and ( id_1674, id_1554, id_1563);
or ( id_1862, id_1853, id_1856, id_1859);
nor ( id_1866, id_1853, id_1856, id_1859);
or ( id_1874, id_1871, id_1872, id_1873);
or ( id_1924, id_1921, id_1922, id_1923);
or ( id_1963, id_1954, id_1957, id_1960);
nor ( id_1967, id_1954, id_1957, id_1960);
or ( id_1975, id_1972, id_1973, id_1974);
or ( id_2013, id_2004, id_2007, id_2010);
nor ( id_2017, id_2004, id_2007, id_2010);
or ( id_2025, id_2022, id_2023, id_2024);
or ( id_2068, id_2059, id_2062, id_2065);
nor ( id_2072, id_2059, id_2062, id_2065);
or ( id_2080, id_2077, id_2078, id_2079);
or ( id_2132, id_2129, id_2130, id_2131);
or ( id_2173, id_2164, id_2167, id_2170);
nor ( id_2177, id_2164, id_2167, id_2170);
or ( id_2185, id_2182, id_2183, id_2184);
or ( id_2225, id_2216, id_2219, id_2222);
nor ( id_2229, id_2216, id_2219, id_2222);
or ( id_2237, id_2234, id_2235, id_2236);
not ( id_2488, id_2485);
not ( id_2679, id_870);
and ( id_2680, id_956, id_870);
not ( id_2698, id_870);
and ( id_2699, id_956, id_870);
not ( id_2717, id_870);
and ( id_2718, id_956, id_870);
not ( id_2734, id_870);
and ( id_2735, id_956, id_870);
not ( id_2752, id_870);
and ( id_2753, id_956, id_870);
not ( id_2769, id_870);
and ( id_2770, id_956, id_870);
not ( id_2786, id_870);
and ( id_2787, id_956, id_870);
not ( id_2803, id_870);
and ( id_2804, id_956, id_870);
or ( id_359, id_917, id_920, id_923);
nor ( id_1029, id_917, id_920, id_923);
nand ( id_565, id_2970, id_2973);
nand ( id_566, id_2967, id_2974);
nand ( id_569, id_2978, id_2981);
nand ( id_570, id_2975, id_2982);
nand ( id_589, id_3050, id_3053);
nand ( id_590, id_3047, id_3054);
nand ( id_595, id_3058, id_3061);
nand ( id_596, id_3055, id_3062);
and ( id_929, id_650, id_926);
and ( id_938, id_630, id_928);
and ( id_944, id_645, id_941);
or ( id_986, id_983, id_984, id_985);
or ( id_1014, id_1011, id_1012, id_1013);
and ( id_1616, id_442, id_1611);
and ( id_1625, id_456, id_1620);
and ( id_1634, id_463, id_1629);
and ( id_1643, id_479, id_1638);
not ( id_360, id_1029);
nand ( id_567, id_565, id_566);
nand ( id_571, id_569, id_570);
buf ( id_579, id_576);
nand ( id_591, id_589, id_590);
nand ( id_597, id_595, id_596);
and ( id_614, id_576, id_610);
not ( id_1240, id_1075);
not ( id_1241, id_1087);
not ( id_1242, id_1099);
not ( id_1243, id_1111);
not ( id_1244, id_1123);
not ( id_1245, id_1135);
not ( id_1246, id_1147);
not ( id_1247, id_1159);
not ( id_1257, id_1075);
not ( id_1258, id_1087);
not ( id_1259, id_1099);
not ( id_1260, id_1111);
not ( id_1261, id_1123);
not ( id_1262, id_1135);
not ( id_1263, id_1147);
not ( id_1264, id_1159);
not ( id_1274, id_1075);
not ( id_1275, id_1087);
not ( id_1276, id_1099);
not ( id_1277, id_1111);
not ( id_1278, id_1123);
not ( id_1279, id_1135);
not ( id_1280, id_1147);
not ( id_1281, id_1159);
not ( id_1291, id_1075);
not ( id_1292, id_1087);
not ( id_1293, id_1099);
not ( id_1294, id_1111);
not ( id_1295, id_1123);
not ( id_1296, id_1135);
not ( id_1297, id_1147);
not ( id_1298, id_1159);
not ( id_1308, id_1075);
not ( id_1309, id_1087);
not ( id_1310, id_1099);
not ( id_1311, id_1111);
not ( id_1312, id_1123);
not ( id_1313, id_1135);
not ( id_1314, id_1147);
not ( id_1315, id_1159);
not ( id_1325, id_1075);
not ( id_1326, id_1087);
not ( id_1327, id_1099);
not ( id_1328, id_1111);
not ( id_1329, id_1123);
not ( id_1330, id_1135);
not ( id_1331, id_1147);
not ( id_1332, id_1159);
not ( id_1342, id_1075);
not ( id_1343, id_1087);
not ( id_1344, id_1099);
not ( id_1345, id_1111);
not ( id_1346, id_1123);
not ( id_1347, id_1135);
not ( id_1348, id_1147);
not ( id_1349, id_1159);
not ( id_1359, id_1075);
not ( id_1360, id_1087);
not ( id_1361, id_1099);
not ( id_1362, id_1111);
not ( id_1363, id_1123);
not ( id_1364, id_1135);
not ( id_1365, id_1147);
not ( id_1366, id_1159);
not ( id_1376, id_1168);
not ( id_1377, id_1177);
not ( id_1378, id_1186);
not ( id_1379, id_1195);
not ( id_1380, id_1204);
not ( id_1381, id_1213);
not ( id_1382, id_1222);
not ( id_1383, id_1231);
not ( id_1393, id_1168);
not ( id_1394, id_1177);
not ( id_1395, id_1186);
not ( id_1396, id_1195);
not ( id_1397, id_1204);
not ( id_1398, id_1213);
not ( id_1399, id_1222);
not ( id_1400, id_1231);
not ( id_1410, id_1168);
not ( id_1411, id_1177);
not ( id_1412, id_1186);
not ( id_1413, id_1195);
not ( id_1414, id_1204);
not ( id_1415, id_1213);
not ( id_1416, id_1222);
not ( id_1417, id_1231);
not ( id_1427, id_1168);
not ( id_1428, id_1177);
not ( id_1429, id_1186);
not ( id_1430, id_1195);
not ( id_1431, id_1204);
not ( id_1432, id_1213);
not ( id_1433, id_1222);
not ( id_1434, id_1231);
not ( id_1444, id_1168);
not ( id_1445, id_1177);
not ( id_1446, id_1186);
not ( id_1447, id_1195);
not ( id_1448, id_1204);
not ( id_1449, id_1213);
not ( id_1450, id_1222);
not ( id_1451, id_1231);
not ( id_1461, id_1168);
not ( id_1462, id_1177);
not ( id_1463, id_1186);
not ( id_1464, id_1195);
not ( id_1465, id_1204);
not ( id_1466, id_1213);
not ( id_1467, id_1222);
not ( id_1468, id_1231);
not ( id_1478, id_1168);
not ( id_1479, id_1177);
not ( id_1480, id_1186);
not ( id_1481, id_1195);
not ( id_1482, id_1204);
not ( id_1483, id_1213);
not ( id_1484, id_1222);
not ( id_1485, id_1231);
not ( id_1495, id_1168);
not ( id_1496, id_1177);
not ( id_1497, id_1186);
not ( id_1498, id_1195);
not ( id_1499, id_1204);
not ( id_1500, id_1213);
not ( id_1501, id_1222);
not ( id_1502, id_1231);
buf ( id_1877, id_1874);
not ( id_1880, id_1874);
not ( id_1891, id_1866);
and ( id_1903, id_986, id_1901);
buf ( id_1927, id_1924);
not ( id_1930, id_1924);
buf ( id_1978, id_1975);
not ( id_1981, id_1975);
not ( id_1992, id_1967);
buf ( id_2028, id_2025);
not ( id_2031, id_2025);
not ( id_2042, id_2017);
buf ( id_2085, id_2080);
not ( id_2088, id_2080);
not ( id_2099, id_2072);
and ( id_2111, id_1014, id_2109);
buf ( id_2137, id_2132);
not ( id_2140, id_2132);
buf ( id_2190, id_2185);
not ( id_2193, id_2185);
not ( id_2204, id_2177);
buf ( id_2242, id_2237);
not ( id_2245, id_2237);
not ( id_2256, id_2229);
and ( id_2320, id_2285, id_1862);
and ( id_2341, id_2289, id_1963);
and ( id_2354, id_2289, id_2013);
and ( id_2367, id_2289, id_2068);
and ( id_2383, id_2298, id_2173);
and ( id_2391, id_2298, id_2225);
not ( id_2474, id_2080);
not ( id_2475, id_2132);
not ( id_2476, id_2185);
not ( id_2477, id_2237);
and ( id_2482, id_2080, id_2132, id_2185, id_2237, id_2481);
nand ( id_361, id_359, id_360);
not ( id_568, id_567);
or ( id_618, id_614, id_616, id_617);
and ( id_1248, id_124, id_1240);
and ( id_1249, id_159, id_1241);
and ( id_1250, id_150, id_1242);
and ( id_1251, id_143, id_1243);
and ( id_1252, id_137, id_1244);
and ( id_1253, id_132, id_1245);
and ( id_1254, id_128, id_1246);
and ( id_1255, id_125, id_1247);
and ( id_1265, id_125, id_1257);
and ( id_1266, id_432, id_1258);
and ( id_1267, id_159, id_1259);
and ( id_1268, id_150, id_1260);
and ( id_1269, id_143, id_1261);
and ( id_1270, id_137, id_1262);
and ( id_1271, id_132, id_1263);
and ( id_1272, id_128, id_1264);
and ( id_1282, id_128, id_1274);
and ( id_1283, id_447, id_1275);
and ( id_1284, id_432, id_1276);
and ( id_1285, id_159, id_1277);
and ( id_1286, id_150, id_1278);
and ( id_1287, id_143, id_1279);
and ( id_1288, id_137, id_1280);
and ( id_1289, id_132, id_1281);
and ( id_1299, id_132, id_1291);
and ( id_1300, id_467, id_1292);
and ( id_1301, id_447, id_1293);
and ( id_1302, id_432, id_1294);
and ( id_1303, id_159, id_1295);
and ( id_1304, id_150, id_1296);
and ( id_1305, id_143, id_1297);
and ( id_1306, id_137, id_1298);
and ( id_1316, id_137, id_1308);
and ( id_1317, id_483, id_1309);
and ( id_1318, id_467, id_1310);
and ( id_1319, id_447, id_1311);
and ( id_1320, id_432, id_1312);
and ( id_1321, id_159, id_1313);
and ( id_1322, id_150, id_1314);
and ( id_1323, id_143, id_1315);
and ( id_1333, id_143, id_1325);
and ( id_1334, id_492, id_1326);
and ( id_1335, id_483, id_1327);
and ( id_1336, id_467, id_1328);
and ( id_1337, id_447, id_1329);
and ( id_1338, id_432, id_1330);
and ( id_1339, id_159, id_1331);
and ( id_1340, id_150, id_1332);
and ( id_1350, id_150, id_1342);
and ( id_1351, id_504, id_1343);
and ( id_1352, id_492, id_1344);
and ( id_1353, id_483, id_1345);
and ( id_1354, id_467, id_1346);
and ( id_1355, id_447, id_1347);
and ( id_1356, id_432, id_1348);
and ( id_1357, id_159, id_1349);
and ( id_1367, id_159, id_1359);
and ( id_1368, id_517, id_1360);
and ( id_1369, id_504, id_1361);
and ( id_1370, id_492, id_1362);
and ( id_1371, id_483, id_1363);
and ( id_1372, id_467, id_1364);
and ( id_1373, id_447, id_1365);
and ( id_1374, id_432, id_1366);
and ( id_1384, id_283, id_1376);
and ( id_1385, id_447, id_1377);
and ( id_1386, id_467, id_1378);
and ( id_1387, id_483, id_1379);
and ( id_1388, id_492, id_1380);
and ( id_1389, id_504, id_1381);
and ( id_1390, id_517, id_1382);
and ( id_1391, id_530, id_1383);
and ( id_1401, id_294, id_1393);
and ( id_1402, id_467, id_1394);
and ( id_1403, id_483, id_1395);
and ( id_1404, id_492, id_1396);
and ( id_1405, id_504, id_1397);
and ( id_1406, id_517, id_1398);
and ( id_1407, id_530, id_1399);
and ( id_1408, id_283, id_1400);
and ( id_1418, id_303, id_1410);
and ( id_1419, id_483, id_1411);
and ( id_1420, id_492, id_1412);
and ( id_1421, id_504, id_1413);
and ( id_1422, id_517, id_1414);
and ( id_1423, id_530, id_1415);
and ( id_1424, id_283, id_1416);
and ( id_1425, id_294, id_1417);
and ( id_1435, id_311, id_1427);
and ( id_1436, id_492, id_1428);
and ( id_1437, id_504, id_1429);
and ( id_1438, id_517, id_1430);
and ( id_1439, id_530, id_1431);
and ( id_1440, id_283, id_1432);
and ( id_1441, id_294, id_1433);
and ( id_1442, id_303, id_1434);
and ( id_1452, id_317, id_1444);
and ( id_1453, id_504, id_1445);
and ( id_1454, id_517, id_1446);
and ( id_1455, id_530, id_1447);
and ( id_1456, id_283, id_1448);
and ( id_1457, id_294, id_1449);
and ( id_1458, id_303, id_1450);
and ( id_1459, id_311, id_1451);
and ( id_1469, id_322, id_1461);
and ( id_1470, id_517, id_1462);
and ( id_1471, id_530, id_1463);
and ( id_1472, id_283, id_1464);
and ( id_1473, id_294, id_1465);
and ( id_1474, id_303, id_1466);
and ( id_1475, id_311, id_1467);
and ( id_1476, id_317, id_1468);
and ( id_1486, id_326, id_1478);
and ( id_1487, id_530, id_1479);
and ( id_1488, id_283, id_1480);
and ( id_1489, id_294, id_1481);
and ( id_1490, id_303, id_1482);
and ( id_1491, id_311, id_1483);
and ( id_1492, id_317, id_1484);
and ( id_1493, id_322, id_1485);
and ( id_1503, id_329, id_1495);
and ( id_1504, id_283, id_1496);
and ( id_1505, id_294, id_1497);
and ( id_1506, id_303, id_1498);
and ( id_1507, id_311, id_1499);
and ( id_1508, id_317, id_1500);
and ( id_1509, id_322, id_1501);
and ( id_1510, id_326, id_1502);
and ( id_2483, id_2474, id_2475, id_2476, id_2477, id_2478);
buf ( id_600, id_597);
and ( id_661, id_568, id_660);
and ( id_669, id_597, id_665);
and ( id_679, id_591, id_678);
nor ( id_1256, id_1248, id_1249, id_1250, id_1251, id_1252, id_1253, id_1254, id_1255);
nor ( id_1273, id_1265, id_1266, id_1267, id_1268, id_1269, id_1270, id_1271, id_1272);
nor ( id_1290, id_1282, id_1283, id_1284, id_1285, id_1286, id_1287, id_1288, id_1289);
nor ( id_1307, id_1299, id_1300, id_1301, id_1302, id_1303, id_1304, id_1305, id_1306);
nor ( id_1324, id_1316, id_1317, id_1318, id_1319, id_1320, id_1321, id_1322, id_1323);
nor ( id_1341, id_1333, id_1334, id_1335, id_1336, id_1337, id_1338, id_1339, id_1340);
nor ( id_1358, id_1350, id_1351, id_1352, id_1353, id_1354, id_1355, id_1356, id_1357);
nor ( id_1375, id_1367, id_1368, id_1369, id_1370, id_1371, id_1372, id_1373, id_1374);
nor ( id_1392, id_1384, id_1385, id_1386, id_1387, id_1388, id_1389, id_1390, id_1391);
nor ( id_1409, id_1401, id_1402, id_1403, id_1404, id_1405, id_1406, id_1407, id_1408);
nor ( id_1426, id_1418, id_1419, id_1420, id_1421, id_1422, id_1423, id_1424, id_1425);
nor ( id_1443, id_1435, id_1436, id_1437, id_1438, id_1439, id_1440, id_1441, id_1442);
nor ( id_1460, id_1452, id_1453, id_1454, id_1455, id_1456, id_1457, id_1458, id_1459);
nor ( id_1477, id_1469, id_1470, id_1471, id_1472, id_1473, id_1474, id_1475, id_1476);
nor ( id_1494, id_1486, id_1487, id_1488, id_1489, id_1490, id_1491, id_1492, id_1493);
nor ( id_1511, id_1503, id_1504, id_1505, id_1506, id_1507, id_1508, id_1509, id_1510);
and ( id_1652, id_618, id_1647);
and ( id_1883, id_169, id_1862, id_1877);
and ( id_1886, id_179, id_1862, id_1880);
and ( id_1889, id_190, id_1866, id_1880);
and ( id_1890, id_200, id_1866, id_1877);
or ( id_1912, id_1903, id_1906, id_1909);
nor ( id_1916, id_1903, id_1906, id_1909);
and ( id_1984, id_169, id_1963, id_1978);
and ( id_1987, id_179, id_1963, id_1981);
and ( id_1990, id_190, id_1967, id_1981);
and ( id_1991, id_200, id_1967, id_1978);
and ( id_2034, id_169, id_2013, id_2028);
and ( id_2037, id_179, id_2013, id_2031);
and ( id_2040, id_190, id_2017, id_2031);
and ( id_2041, id_200, id_2017, id_2028);
and ( id_2091, id_169, id_2068, id_2085);
and ( id_2094, id_179, id_2068, id_2088);
and ( id_2097, id_190, id_2072, id_2088);
and ( id_2098, id_200, id_2072, id_2085);
or ( id_2120, id_2111, id_2114, id_2117);
nor ( id_2124, id_2111, id_2114, id_2117);
and ( id_2196, id_169, id_2173, id_2190);
and ( id_2199, id_179, id_2173, id_2193);
and ( id_2202, id_190, id_2177, id_2193);
and ( id_2203, id_200, id_2177, id_2190);
and ( id_2248, id_169, id_2225, id_2242);
and ( id_2251, id_179, id_2225, id_2245);
and ( id_2254, id_190, id_2229, id_2245);
and ( id_2255, id_200, id_2229, id_2242);
or ( id_2484, id_2482, id_2483);
buf ( id_2991, id_571);
buf ( id_2994, id_579);
buf ( id_2999, id_571);
buf ( id_3002, id_579);
buf ( id_3063, id_591);
buf ( id_3071, id_591);
buf ( id_3124, id_2320);
buf ( id_3134, id_2320);
buf ( id_3158, id_2341);
buf ( id_3166, id_2341);
buf ( id_3174, id_2354);
buf ( id_3182, id_2354);
buf ( id_3190, id_2367);
buf ( id_3200, id_2367);
buf ( id_3224, id_2383);
buf ( id_3232, id_2383);
buf ( id_3240, id_2391);
buf ( id_3248, id_2391);
nor ( id_663, id_661, id_662);
or ( id_673, id_669, id_671, id_672);
nor ( id_681, id_679, id_680);
and ( id_1536, id_1256, id_1533);
and ( id_1537, id_1392, id_1534);
and ( id_1582, id_1273, id_1581);
and ( id_1583, id_1409, id_1512);
and ( id_1586, id_1290, id_1585);
and ( id_1587, id_1426, id_1512);
and ( id_1590, id_1307, id_1589);
and ( id_1591, id_1443, id_1512);
and ( id_1594, id_1324, id_1593);
and ( id_1595, id_1460, id_1512);
and ( id_1598, id_1341, id_1597);
and ( id_1599, id_1477, id_1512);
and ( id_1602, id_1358, id_1601);
and ( id_1603, id_1494, id_1512);
and ( id_1606, id_1375, id_1605);
and ( id_1607, id_1511, id_1512);
or ( id_1894, id_1889, id_1890, id_1891);
or ( id_1997, id_1990, id_1991, id_1992);
or ( id_2047, id_2040, id_2041, id_2042);
or ( id_2102, id_2097, id_2098, id_2099);
or ( id_2209, id_2202, id_2203, id_2204);
or ( id_2261, id_2254, id_2255, id_2256);
and ( id_2489, id_2484, id_2488);
not ( id_3005, id_2999);
not ( id_3006, id_3002);
not ( id_3077, id_3071);
not ( id_3069, id_3063);
not ( id_2997, id_2991);
not ( id_2998, id_2994);
and ( id_689, id_681, id_683);
and ( id_700, id_663, id_694);
or ( id_1539, id_1536, id_1537, id_1538);
or ( id_1584, id_1582, id_1583);
or ( id_1588, id_1586, id_1587);
or ( id_1592, id_1590, id_1591);
or ( id_1596, id_1594, id_1595);
or ( id_1600, id_1598, id_1599);
or ( id_1604, id_1602, id_1603);
or ( id_1608, id_1606, id_1607);
and ( id_1661, id_673, id_1656);
or ( id_1892, id_1883, id_1886);
nor ( id_1893, id_1883, id_1886);
and ( id_1933, id_169, id_1912, id_1927);
and ( id_1936, id_179, id_1912, id_1930);
and ( id_1939, id_190, id_1916, id_1930);
and ( id_1940, id_200, id_1916, id_1927);
not ( id_1941, id_1916);
or ( id_1993, id_1984, id_1987);
nor ( id_1996, id_1984, id_1987);
or ( id_2043, id_2034, id_2037);
nor ( id_2046, id_2034, id_2037);
or ( id_2100, id_2091, id_2094);
nor ( id_2101, id_2091, id_2094);
and ( id_2143, id_169, id_2120, id_2137);
and ( id_2146, id_179, id_2120, id_2140);
and ( id_2149, id_190, id_2124, id_2140);
and ( id_2150, id_200, id_2124, id_2137);
not ( id_2151, id_2124);
or ( id_2205, id_2196, id_2199);
nor ( id_2208, id_2196, id_2199);
or ( id_2257, id_2248, id_2251);
nor ( id_2260, id_2248, id_2251);
not ( id_3138, id_3134);
and ( id_2328, id_2285, id_1912);
not ( id_3162, id_3158);
not ( id_3170, id_3166);
not ( id_3178, id_3174);
not ( id_3186, id_3182);
not ( id_3204, id_3200);
and ( id_2375, id_2298, id_2120);
not ( id_3236, id_3232);
not ( id_3244, id_3240);
not ( id_3252, id_3248);
not ( id_3228, id_3224);
buf ( id_3066, id_600);
buf ( id_3074, id_600);
not ( id_3128, id_3124);
not ( id_3194, id_3190);
nand ( id_619, id_2994, id_2997);
nand ( id_620, id_2991, id_2998);
nand ( id_582, id_3002, id_3005);
nand ( id_583, id_2999, id_3006);
or ( id_692, id_689, id_690, id_691);
or ( id_703, id_700, id_701, id_702);
and ( id_1612, id_1539, id_1609);
and ( id_1621, id_1584, id_1618);
and ( id_1630, id_1588, id_1627);
and ( id_1639, id_1592, id_1636);
and ( id_1648, id_1596, id_1645);
and ( id_1657, id_1600, id_1654);
and ( id_1666, id_1604, id_1663);
and ( id_1675, id_1608, id_1672);
and ( id_1895, id_1893, id_1894);
or ( id_1946, id_1939, id_1940, id_1941);
and ( id_1998, id_1996, id_1997);
and ( id_2048, id_2046, id_2047);
and ( id_2103, id_2101, id_2102);
or ( id_2156, id_2149, id_2150, id_2151);
and ( id_2210, id_2208, id_2209);
and ( id_2262, id_2260, id_2261);
not ( id_2271, id_1892);
not ( id_2311, id_2100);
nand ( id_356, id_619, id_620);
nand ( id_357, id_582, id_583);
nand ( id_603, id_3074, id_3077);
not ( id_3078, id_3074);
nand ( id_606, id_3066, id_3069);
not ( id_3070, id_3066);
and ( id_1670, id_703, id_1665);
and ( id_1679, id_692, id_1674);
or ( id_1942, id_1933, id_1936);
nor ( id_1945, id_1933, id_1936);
or ( id_2152, id_2143, id_2146);
nor ( id_2155, id_2143, id_2146);
and ( id_2445, id_1993, id_2293);
and ( id_2448, id_2043, id_2293);
and ( id_2455, id_2205, id_2302);
and ( id_2458, id_2257, id_2302);
buf ( id_3142, id_2328);
buf ( id_3150, id_2328);
buf ( id_3208, id_2375);
buf ( id_3216, id_2375);
nand ( id_358, id_356, id_357);
nand ( id_604, id_3071, id_3078);
nand ( id_607, id_3063, id_3070);
and ( id_1947, id_1945, id_1946);
and ( id_2157, id_2155, id_2156);
buf ( id_2317, id_1895);
buf ( id_2338, id_1998);
buf ( id_2351, id_2048);
buf ( id_2364, id_2103);
buf ( id_2380, id_2210);
buf ( id_2388, id_2262);
nand ( id_605, id_603, id_604);
nand ( id_608, id_606, id_607);
nand ( id_2272, id_1895, id_1942);
nand ( id_2312, id_2103, id_2152);
not ( id_3146, id_3142);
not ( id_3154, id_3150);
not ( id_3220, id_3216);
not ( id_3212, id_3208);
and ( id_2444, id_1942, id_2288);
buf ( id_2451, id_2448);
and ( id_2454, id_2152, id_2293);
buf ( id_2461, id_2458);
not ( id_2530, id_2445);
buf ( id_3323, id_2458);
not ( id_349, id_605);
not ( id_350, id_608);
and ( id_2265, id_1895, id_1947, id_1998, id_2048);
nand ( id_2273, id_1895, id_1947, id_1993);
nand ( id_2274, id_2043, id_1947, id_1998, id_1895);
and ( id_2309, id_2103, id_2157, id_2210, id_2262);
nand ( id_2313, id_2103, id_2157, id_2205);
nand ( id_2314, id_2257, id_2157, id_2210, id_2103);
buf ( id_2325, id_1947);
buf ( id_2372, id_2157);
not ( id_2523, id_2444);
not ( id_2533, id_2454);
buf ( id_3121, id_2317);
buf ( id_3131, id_2317);
buf ( id_3155, id_2338);
buf ( id_3163, id_2338);
buf ( id_3171, id_2351);
buf ( id_3179, id_2351);
buf ( id_3187, id_2364);
buf ( id_3197, id_2364);
buf ( id_3221, id_2380);
buf ( id_3229, id_2380);
buf ( id_3237, id_2388);
buf ( id_3245, id_2388);
nand ( id_351, id_349, id_350);
nand ( id_2275, id_2271, id_2272, id_2273, id_2274);
nand ( id_2315, id_2311, id_2312, id_2313, id_2314);
not ( id_3329, id_3323);
and ( id_372, id_2309, id_2265);
nand ( id_2324, id_3131, id_3138);
nand ( id_2350, id_3163, id_3170);
nand ( id_2363, id_3179, id_3186);
nand ( id_2371, id_3197, id_3204);
nand ( id_2387, id_3229, id_3236);
nand ( id_2400, id_3245, id_3252);
buf ( id_2268, id_2265);
not ( id_3137, id_3131);
not ( id_3161, id_3155);
nand ( id_2345, id_3155, id_3162);
not ( id_3169, id_3163);
not ( id_3177, id_3171);
nand ( id_2358, id_3171, id_3178);
not ( id_3185, id_3179);
not ( id_3203, id_3197);
not ( id_3235, id_3229);
not ( id_3243, id_3237);
nand ( id_2395, id_3237, id_3244);
not ( id_3251, id_3245);
not ( id_3227, id_3221);
nand ( id_2432, id_3221, id_3228);
and ( id_2490, id_2309, id_2485);
not ( id_3127, id_3121);
nand ( id_3130, id_3121, id_3128);
buf ( id_3139, id_2325);
buf ( id_3147, id_2325);
not ( id_3193, id_3187);
nand ( id_3196, id_3187, id_3194);
buf ( id_3205, id_2372);
buf ( id_3213, id_2372);
nand ( id_2307, id_2265, id_2315);
not ( id_2308, id_2275);
nand ( id_2323, id_3134, id_3137);
nand ( id_2349, id_3166, id_3169);
nand ( id_2362, id_3182, id_3185);
nand ( id_2370, id_3200, id_3203);
nand ( id_2386, id_3232, id_3235);
nand ( id_2399, id_3248, id_3251);
nand ( id_2344, id_3158, id_3161);
nand ( id_2357, id_3174, id_3177);
nand ( id_2394, id_3240, id_3243);
nand ( id_2431, id_3224, id_3227);
and ( id_2464, id_2315, id_2302);
or ( id_2491, id_2489, id_2490);
nand ( id_3129, id_3124, id_3127);
nand ( id_3195, id_3190, id_3193);
and ( id_368, id_2307, id_2308);
nand ( id_1615, id_2323, id_2324);
nand ( id_2337, id_3147, id_3154);
nand ( id_1633, id_2349, id_2350);
nand ( id_1642, id_2362, id_2363);
nand ( id_1651, id_2370, id_2371);
nand ( id_2379, id_3213, id_3220);
nand ( id_1669, id_2386, id_2387);
nand ( id_1678, id_2399, id_2400);
not ( id_3145, id_3139);
nand ( id_2332, id_3139, id_3146);
not ( id_3153, id_3147);
nand ( id_2346, id_2344, id_2345);
nand ( id_2359, id_2357, id_2358);
not ( id_3219, id_3213);
nand ( id_2396, id_2394, id_2395);
not ( id_3211, id_3205);
nand ( id_2425, id_3205, id_3212);
nand ( id_2433, id_2431, id_2432);
nand ( id_3272, id_3129, id_3130);
nand ( id_3308, id_3195, id_3196);
not ( id_369, id_368);
not ( id_1613, id_1615);
nand ( id_2336, id_3150, id_3153);
not ( id_1631, id_1633);
not ( id_1640, id_1642);
not ( id_1649, id_1651);
nand ( id_2378, id_3216, id_3219);
not ( id_1667, id_1669);
not ( id_1676, id_1678);
nand ( id_2331, id_3142, id_3145);
nand ( id_2424, id_3208, id_3211);
buf ( id_2467, id_2464);
buf ( id_2495, id_2491);
buf ( id_3295, id_2464);
and ( id_3374, id_330, id_2491);
and ( id_1614, id_1613, id_1610);
nand ( id_1624, id_2336, id_2337);
and ( id_1632, id_1631, id_1628);
and ( id_1641, id_1640, id_1637);
and ( id_1650, id_1649, id_1646);
nand ( id_1660, id_2378, id_2379);
and ( id_1668, id_1667, id_1664);
and ( id_1677, id_1676, id_1673);
nand ( id_2333, id_2331, id_2332);
buf ( id_2406, id_2346);
buf ( id_2409, id_2346);
buf ( id_2415, id_2359);
buf ( id_2419, id_2359);
nand ( id_2426, id_2424, id_2425);
buf ( id_2439, id_2396);
and ( id_2518, id_2433, id_2461);
not ( id_3276, id_3272);
not ( id_3312, id_3308);
and ( id_2612, id_330, id_2396);
buf ( id_3326, id_2433);
nor ( id_1617, id_1612, id_1614, id_1616);
not ( id_1622, id_1624);
nor ( id_1635, id_1630, id_1632, id_1634);
nor ( id_1644, id_1639, id_1641, id_1643);
nor ( id_1653, id_1648, id_1650, id_1652);
not ( id_1658, id_1660);
nor ( id_1671, id_1666, id_1668, id_1670);
nor ( id_1680, id_1675, id_1677, id_1679);
and ( id_2500, id_2467, id_2268);
and ( id_2505, id_2495, id_2268);
or ( id_2519, id_2455, id_2518);
not ( id_3378, id_3374);
not ( id_2642, id_2467);
buf ( id_2645, id_2467);
not ( id_3301, id_3295);
and ( id_1623, id_1622, id_1619);
and ( id_1659, id_1658, id_1655);
buf ( id_2401, id_2333);
or ( id_2501, id_2275, id_2500);
and ( id_2511, id_2495, id_2419, id_2409);
and ( id_2512, id_2495, id_2415);
and ( id_2513, id_2439, id_2433, id_2426);
and ( id_2514, id_2439, id_2433);
and ( id_2517, id_2467, id_2415);
nand ( id_2531, id_2409, id_2451);
nand ( id_2532, id_2409, id_2419, id_2467);
nand ( id_2534, id_2426, id_2455);
nand ( id_2535, id_2426, id_2433, id_2461);
nand ( id_2607, id_3326, id_3329);
not ( id_3330, id_3326);
and ( id_2643, id_330, id_2491, id_2642);
and ( id_2687, id_1617, id_2680);
and ( id_2725, id_1635, id_2718);
and ( id_2742, id_1644, id_2735);
and ( id_2760, id_1653, id_2753);
and ( id_2794, id_1671, id_2787);
and ( id_2811, id_1680, id_2804);
buf ( id_3280, id_2333);
buf ( id_3290, id_2409);
buf ( id_3298, id_2415);
buf ( id_3316, id_2426);
buf ( id_3406, id_2612);
buf ( id_3414, id_2612);
and ( id_3422, id_2439, id_2439);
nor ( id_1626, id_1621, id_1623, id_1625);
nor ( id_1662, id_1657, id_1659, id_1661);
and ( id_2567, id_330, id_2512);
and ( id_2589, id_330, id_2513);
nand ( id_2608, id_3323, id_3330);
buf ( id_2654, id_2519);
buf ( id_3253, id_2505);
nand ( id_3277, id_2530, id_2531, id_2532);
or ( id_3287, id_2448, id_2517);
nand ( id_3305, id_2533, id_2534, id_2535);
buf ( id_3313, id_2519);
and ( id_3350, id_330, id_2511);
or ( id_932, id_2643, id_2645);
and ( id_2508, id_2495, id_2401, id_2409, id_2419);
nand ( id_2524, id_2401, id_2445);
nand ( id_2525, id_2401, id_2406, id_2451);
nand ( id_2526, id_2401, id_2406, id_2419, id_2467);
not ( id_3294, id_3290);
nand ( id_2609, id_2607, id_2608);
not ( id_3410, id_3406);
not ( id_3418, id_3414);
nand ( id_2624, id_3422, id_3425);
not ( id_3426, id_3422);
buf ( id_2629, id_2501);
nor ( id_2647, id_2643, id_2645);
and ( id_2706, id_1626, id_2699);
and ( id_2777, id_1662, id_2770);
buf ( id_3264, id_2501);
not ( id_3284, id_3280);
not ( id_3302, id_3298);
nand ( id_3303, id_3298, id_3301);
not ( id_3320, id_3316);
and ( id_3398, id_330, id_2514);
not ( id_2657, id_2654);
and ( id_398, id_2519, id_2654);
and ( id_933, id_932, id_927);
nand ( id_2527, id_2523, id_2524, id_2525, id_2526);
not ( id_3259, id_3253);
not ( id_3354, id_3350);
not ( id_3293, id_3287);
nand ( id_2563, id_3287, id_3294);
not ( id_3311, id_3305);
nand ( id_2585, id_3305, id_3312);
nand ( id_2625, id_3419, id_3426);
not ( id_3283, id_3277);
nand ( id_3286, id_3277, id_3284);
nand ( id_3304, id_3295, id_3302);
not ( id_3319, id_3313);
nand ( id_3322, id_3313, id_3320);
buf ( id_3358, id_2567);
buf ( id_3366, id_2567);
buf ( id_3382, id_2589);
buf ( id_3390, id_2589);
and ( id_397, id_330, id_2514, id_2657);
and ( id_2544, id_330, id_2508);
nand ( id_2562, id_3290, id_3293);
nand ( id_2584, id_3308, id_3311);
not ( id_3402, id_3398);
nand ( id_2626, id_2624, id_2625);
not ( id_2632, id_2629);
and ( id_2634, id_2501, id_2629);
buf ( id_2650, id_2647);
not ( id_3268, id_3264);
buf ( id_3256, id_2508);
nand ( id_3285, id_3280, id_3283);
nand ( id_3321, id_3316, id_3319);
nand ( id_3371, id_3303, id_3304);
buf ( id_3403, id_2609);
buf ( id_3411, id_2609);
or ( id_362, id_929, id_933, id_938);
nor ( id_1030, id_929, id_933, id_938);
or ( id_399, id_397, id_398);
nand ( id_2564, id_2562, id_2563);
not ( id_3362, id_3358);
not ( id_3370, id_3366);
nand ( id_2586, id_2584, id_2585);
not ( id_3386, id_3382);
not ( id_3394, id_3390);
and ( id_2633, id_330, id_2505, id_2632);
buf ( id_3261, id_2527);
buf ( id_3269, id_2527);
nand ( id_3347, id_3285, id_3286);
nand ( id_3395, id_3321, id_3322);
not ( id_363, id_1030);
nand ( id_2536, id_3256, id_3259);
not ( id_3260, id_3256);
not ( id_3377, id_3371);
nand ( id_2580, id_3371, id_3378);
not ( id_3409, id_3403);
nand ( id_2616, id_3403, id_3410);
not ( id_3417, id_3411);
nand ( id_2622, id_3411, id_3418);
nor ( id_2635, id_2633, id_2634);
and ( id_2805, id_2626, id_2802);
and ( id_2808, id_2626, id_2803);
buf ( id_3334, id_2544);
buf ( id_3342, id_2544);
buf ( id_3454, id_2650);
and ( id_364, id_362, id_363);
nand ( id_2537, id_3253, id_3260);
not ( id_3275, id_3269);
nand ( id_2540, id_3269, id_3276);
not ( id_3353, id_3347);
nand ( id_2557, id_3347, id_3354);
nand ( id_2579, id_3374, id_3377);
not ( id_3401, id_3395);
nand ( id_2602, id_3395, id_3402);
nand ( id_2615, id_3406, id_3409);
nand ( id_2621, id_3414, id_3417);
not ( id_3267, id_3261);
nand ( id_3112, id_3261, id_3268);
buf ( id_3355, id_2564);
buf ( id_3363, id_2564);
buf ( id_3379, id_2586);
buf ( id_3387, id_2586);
nand ( id_2538, id_2536, id_2537);
nand ( id_2539, id_3272, id_3275);
not ( id_3338, id_3334);
not ( id_3346, id_3342);
nand ( id_2556, id_3350, id_3353);
nand ( id_2581, id_2579, id_2580);
nand ( id_2601, id_3398, id_3401);
nand ( id_2617, id_2615, id_2616);
nand ( id_2623, id_2621, id_2622);
buf ( id_2638, id_2635);
not ( id_3458, id_3454);
or ( id_2814, id_2805, id_2808, id_2811);
nor ( id_2816, id_2805, id_2808, id_2811);
nand ( id_3111, id_3264, id_3267);
nand ( id_2541, id_2539, id_2540);
nand ( id_2558, id_2556, id_2557);
not ( id_3361, id_3355);
nand ( id_2571, id_3355, id_3362);
not ( id_3369, id_3363);
nand ( id_2577, id_3363, id_3370);
not ( id_3385, id_3379);
nand ( id_2593, id_3379, id_3386);
not ( id_3393, id_3387);
nand ( id_2598, id_3387, id_3394);
nand ( id_2603, id_2601, id_2602);
nand ( id_3113, id_3111, id_3112);
and ( id_3116, id_330, id_2538);
not ( id_3451, id_2623);
not ( id_395, id_2816);
nand ( id_2570, id_3358, id_3361);
nand ( id_2576, id_3366, id_3369);
nand ( id_2592, id_3382, id_3385);
nand ( id_2597, id_3390, id_3393);
and ( id_2736, id_2581, id_2733);
and ( id_2739, id_2581, id_2734);
and ( id_2788, id_2617, id_2785);
buf ( id_3438, id_2638);
and ( id_3446, id_2617, id_2647);
buf ( id_3459, id_2814);
and ( id_396, id_2814, id_395);
not ( id_3119, id_3113);
not ( id_3120, id_3116);
nand ( id_2572, id_2570, id_2571);
nand ( id_2578, id_2576, id_2577);
nand ( id_2594, id_2592, id_2593);
nand ( id_2599, id_2597, id_2598);
nand ( id_2677, id_3451, id_3458);
not ( id_3457, id_3451);
and ( id_2700, id_2558, id_2697);
and ( id_2771, id_2603, id_2768);
buf ( id_3331, id_2541);
buf ( id_3339, id_2541);
buf ( id_3427, id_2558);
buf ( id_3443, id_2603);
nand ( id_954, id_3116, id_3119);
nand ( id_955, id_3113, id_3120);
not ( id_2600, id_2599);
not ( id_3442, id_3438);
not ( id_3450, id_3446);
nand ( id_2676, id_3454, id_3457);
or ( id_2745, id_2736, id_2739, id_2742);
nor ( id_2748, id_2736, id_2739, id_2742);
not ( id_3465, id_3459);
not ( id_3435, id_2578);
nand ( id_950, id_954, id_955);
not ( id_3337, id_3331);
nand ( id_2548, id_3331, id_3338);
not ( id_3345, id_3339);
nand ( id_2553, id_3339, id_3346);
nor ( id_2661, id_2600, id_2650);
and ( id_2662, id_2617, id_2603, id_2594, id_2650);
not ( id_3433, id_3427);
not ( id_3449, id_3443);
nand ( id_2672, id_3443, id_3450);
nand ( id_2674, id_2676, id_2677);
and ( id_2719, id_2572, id_2716);
and ( id_2754, id_2594, id_2751);
and ( id_3430, id_2572, id_2635);
not ( id_383, id_2748);
and ( id_951, id_950, id_943);
nand ( id_2547, id_3334, id_3337);
nand ( id_2552, id_3342, id_3345);
or ( id_2663, id_2661, id_2662);
nand ( id_2670, id_3435, id_3442);
not ( id_3441, id_3435);
nand ( id_2671, id_3446, id_3449);
not ( id_2675, id_2674);
buf ( id_3491, id_2745);
buf ( id_3499, id_2745);
and ( id_384, id_2745, id_383);
nand ( id_2549, id_2547, id_2548);
nand ( id_2554, id_2552, id_2553);
nand ( id_2664, id_3430, id_3433);
not ( id_3434, id_3430);
nand ( id_2669, id_3438, id_3441);
nand ( id_2673, id_2671, id_2672);
and ( id_2757, id_2663, id_2752);
and ( id_2791, id_2675, id_2786);
or ( id_365, id_944, id_947, id_951);
nor ( id_1031, id_944, id_947, id_951);
not ( id_2555, id_2554);
nand ( id_2665, id_3427, id_3434);
nand ( id_2667, id_2669, id_2670);
and ( id_2774, id_2673, id_2769);
not ( id_3497, id_3491);
not ( id_3505, id_3499);
not ( id_366, id_1031);
nor ( id_2658, id_2555, id_2638);
and ( id_2659, id_2572, id_2558, id_2549, id_2638);
nand ( id_2666, id_2664, id_2665);
not ( id_2668, id_2667);
and ( id_2681, id_2549, id_2678);
or ( id_2763, id_2754, id_2757, id_2760);
nor ( id_2765, id_2754, id_2757, id_2760);
or ( id_2797, id_2788, id_2791, id_2794);
nor ( id_2799, id_2788, id_2791, id_2794);
and ( id_367, id_365, id_366);
or ( id_2660, id_2658, id_2659);
and ( id_2703, id_2666, id_2698);
and ( id_2722, id_2668, id_2717);
or ( id_2780, id_2771, id_2774, id_2777);
nor ( id_2782, id_2771, id_2774, id_2777);
not ( id_386, id_2765);
not ( id_392, id_2799);
and ( id_2684, id_2660, id_2679);
buf ( id_3462, id_2797);
buf ( id_3470, id_2763);
and ( id_387, id_2763, id_386);
not ( id_389, id_2782);
and ( id_393, id_2797, id_392);
or ( id_2709, id_2700, id_2703, id_2706);
nor ( id_2713, id_2700, id_2703, id_2706);
or ( id_2728, id_2719, id_2722, id_2725);
nor ( id_2730, id_2719, id_2722, id_2725);
and ( id_2922, id_2816, id_2799, id_2782, id_2765);
buf ( id_3467, id_2780);
and ( id_390, id_2780, id_389);
or ( id_2690, id_2681, id_2684, id_2687);
nor ( id_2694, id_2681, id_2684, id_2687);
nand ( id_2821, id_3462, id_3465);
not ( id_3466, id_3462);
not ( id_3474, id_3470);
and ( id_378, id_2709, id_2709);
not ( id_380, id_2730);
nand ( id_2822, id_3459, id_3466);
not ( id_3473, id_3467);
nand ( id_2827, id_3467, id_3474);
buf ( id_2839, id_2728);
and ( id_2883, id_2709, id_2871);
buf ( id_3507, id_2709);
and ( id_375, id_2690, id_2690);
and ( id_381, id_2728, id_380);
nand ( id_2823, id_2821, id_2822);
nand ( id_2826, id_3470, id_3473);
and ( id_2880, id_2871, id_2690);
and ( id_2925, id_2748, id_2730, id_2713, id_2694);
and ( id_2928, id_2713, id_2694, id_2874);
buf ( id_3510, id_2690);
nand ( id_2828, id_2826, id_2827);
buf ( id_3494, id_2839);
buf ( id_3502, id_2839);
not ( id_3513, id_3507);
buf ( id_3544, id_2883);
buf ( id_3552, id_2883);
and ( id_406, id_2922, id_2925);
and ( id_2929, id_2922, id_2925);
buf ( id_3475, id_2823);
buf ( id_3483, id_2823);
not ( id_3514, id_3510);
nand ( id_3515, id_3510, id_3513);
buf ( id_3541, id_2880);
buf ( id_3549, id_2880);
not ( id_407, id_406);
nor ( id_2930, id_2928, id_2929);
nand ( id_2842, id_3494, id_3497);
not ( id_3498, id_3494);
nand ( id_2852, id_3502, id_3505);
not ( id_3506, id_3502);
not ( id_3548, id_3544);
not ( id_3556, id_3552);
buf ( id_3478, id_2828);
buf ( id_3486, id_2828);
nand ( id_3516, id_3507, id_3514);
and ( id_408, id_213, id_2930);
not ( id_3481, id_3475);
not ( id_3489, id_3483);
nand ( id_2843, id_3491, id_3498);
nand ( id_2853, id_3499, id_3506);
not ( id_3547, id_3541);
nand ( id_2887, id_3541, id_3548);
nand ( id_2896, id_3549, id_3556);
not ( id_3555, id_3549);
nand ( id_3520, id_3515, id_3516);
not ( id_409, id_408);
nand ( id_2831, id_3478, id_3481);
not ( id_3482, id_3478);
nand ( id_2836, id_3486, id_3489);
not ( id_3490, id_3486);
nand ( id_2844, id_2842, id_2843);
nand ( id_2848, id_2852, id_2853);
nand ( id_2886, id_3544, id_3547);
nand ( id_2895, id_3552, id_3555);
nand ( id_2832, id_3475, id_3482);
nand ( id_2837, id_3483, id_3490);
not ( id_2849, id_2848);
not ( id_3524, id_3520);
nand ( id_2888, id_2886, id_2887);
nand ( id_2891, id_2895, id_2896);
nand ( id_2833, id_2831, id_2832);
nand ( id_2838, id_2836, id_2837);
not ( id_2892, id_2891);
buf ( id_3517, id_2844);
and ( id_2906, id_2844, id_2888, id_2900);
and ( id_2908, id_2849, id_2888, id_2903);
not ( id_2913, id_2838);
not ( id_3523, id_3517);
nand ( id_2855, id_3517, id_3524);
and ( id_2907, id_2844, id_2892, id_2903);
and ( id_2909, id_2849, id_2892, id_2900);
buf ( id_3525, id_2833);
buf ( id_3533, id_2833);
nand ( id_2854, id_3520, id_3523);
or ( id_2910, id_2906, id_2907, id_2908, id_2909);
buf ( id_3560, id_2913);
buf ( id_3568, id_2913);
nand ( id_2856, id_2854, id_2855);
not ( id_3539, id_3533);
not ( id_3531, id_3525);
not ( id_3572, id_3568);
not ( id_3564, id_3560);
buf ( id_3557, id_2910);
buf ( id_3565, id_2910);
buf ( id_3528, id_2856);
buf ( id_3536, id_2856);
nand ( id_2921, id_3557, id_3564);
nand ( id_2917, id_3565, id_3572);
not ( id_3571, id_3565);
not ( id_3563, id_3557);
nand ( id_2863, id_3528, id_3531);
nand ( id_2859, id_3536, id_3539);
nand ( id_2920, id_3560, id_3563);
nand ( id_2916, id_3568, id_3571);
not ( id_3540, id_3536);
not ( id_3532, id_3528);
nand ( id_2864, id_3525, id_3532);
nand ( id_2860, id_3533, id_3540);
nand ( id_403, id_2920, id_2921);
nand ( id_404, id_2916, id_2917);
nand ( id_400, id_2863, id_2864);
nand ( id_401, id_2859, id_2860);
and ( id_405, id_403, id_404);
nand ( id_402, id_400, id_401);

endmodule
