module c6288nr
( id_1gat ,id_18gat ,id_35gat ,id_52gat ,id_69gat ,id_86gat ,id_103gat ,id_120gat ,id_137gat ,id_154gat ,id_171gat ,id_188gat ,id_205gat ,id_222gat ,id_239gat ,id_256gat ,id_273gat ,id_290gat ,id_307gat ,id_324gat ,id_341gat ,id_358gat ,id_375gat ,id_392gat ,id_409gat ,id_426gat ,id_443gat ,id_460gat ,id_477gat ,id_494gat ,id_511gat ,id_528gat ,id_545gat ,id_1581gat ,id_1901gat ,id_2223gat ,id_2548gat ,id_2877gat ,id_3211gat ,id_3552gat ,id_3895gat ,id_4241gat ,id_4591gat ,id_4946gat ,id_5308gat ,id_5672gat ,id_5971gat ,id_6123gat ,id_6150gat ,id_6160gat ,id_6170gat ,id_6180gat ,id_6190gat ,id_6200gat ,id_6210gat ,id_6220gat ,id_6230gat ,id_6240gat ,id_6250gat ,id_6260gat ,id_6270gat ,id_6280gat ,id_6287gat ,id_6288gat  );

input id_1gat, id_18gat, id_35gat, id_52gat, id_69gat, id_86gat, id_103gat, id_120gat, id_137gat, id_154gat, id_171gat, id_188gat, id_205gat, id_222gat, id_239gat, id_256gat, id_273gat, id_290gat, id_307gat, id_324gat, id_341gat, id_358gat, id_375gat, id_392gat, id_409gat, id_426gat, id_443gat, id_460gat, id_477gat, id_494gat, id_511gat, id_528gat;

output id_545gat, id_1581gat, id_1901gat, id_2223gat, id_2548gat, id_2877gat, id_3211gat, id_3552gat, id_3895gat, id_4241gat, id_4591gat, id_4946gat, id_5308gat, id_5672gat, id_5971gat, id_6123gat, id_6150gat, id_6160gat, id_6170gat, id_6180gat, id_6190gat, id_6200gat, id_6210gat, id_6220gat, id_6230gat, id_6240gat, id_6250gat, id_6260gat, id_6270gat, id_6280gat, id_6287gat, id_6288gat;

and ( id_545gat, id_1gat, id_273gat);
and ( id_546gat, id_1gat, id_290gat);
and ( id_549gat, id_1gat, id_307gat);
and ( id_552gat, id_1gat, id_324gat);
and ( id_555gat, id_1gat, id_341gat);
and ( id_558gat, id_1gat, id_358gat);
and ( id_561gat, id_1gat, id_375gat);
and ( id_564gat, id_1gat, id_392gat);
and ( id_567gat, id_1gat, id_409gat);
and ( id_570gat, id_1gat, id_426gat);
and ( id_573gat, id_1gat, id_443gat);
and ( id_576gat, id_1gat, id_460gat);
and ( id_579gat, id_1gat, id_477gat);
and ( id_582gat, id_1gat, id_494gat);
and ( id_585gat, id_1gat, id_511gat);
and ( id_588gat, id_1gat, id_528gat);
and ( id_591gat, id_18gat, id_273gat);
and ( id_594gat, id_18gat, id_290gat);
and ( id_597gat, id_18gat, id_307gat);
and ( id_600gat, id_18gat, id_324gat);
and ( id_603gat, id_18gat, id_341gat);
and ( id_606gat, id_18gat, id_358gat);
and ( id_609gat, id_18gat, id_375gat);
and ( id_612gat, id_18gat, id_392gat);
and ( id_615gat, id_18gat, id_409gat);
and ( id_618gat, id_18gat, id_426gat);
and ( id_621gat, id_18gat, id_443gat);
and ( id_624gat, id_18gat, id_460gat);
and ( id_627gat, id_18gat, id_477gat);
and ( id_630gat, id_18gat, id_494gat);
and ( id_633gat, id_18gat, id_511gat);
and ( id_636gat, id_18gat, id_528gat);
and ( id_639gat, id_35gat, id_273gat);
and ( id_642gat, id_35gat, id_290gat);
and ( id_645gat, id_35gat, id_307gat);
and ( id_648gat, id_35gat, id_324gat);
and ( id_651gat, id_35gat, id_341gat);
and ( id_654gat, id_35gat, id_358gat);
and ( id_657gat, id_35gat, id_375gat);
and ( id_660gat, id_35gat, id_392gat);
and ( id_663gat, id_35gat, id_409gat);
and ( id_666gat, id_35gat, id_426gat);
and ( id_669gat, id_35gat, id_443gat);
and ( id_672gat, id_35gat, id_460gat);
and ( id_675gat, id_35gat, id_477gat);
and ( id_678gat, id_35gat, id_494gat);
and ( id_681gat, id_35gat, id_511gat);
and ( id_684gat, id_35gat, id_528gat);
and ( id_687gat, id_52gat, id_273gat);
and ( id_690gat, id_52gat, id_290gat);
and ( id_693gat, id_52gat, id_307gat);
and ( id_696gat, id_52gat, id_324gat);
and ( id_699gat, id_52gat, id_341gat);
and ( id_702gat, id_52gat, id_358gat);
and ( id_705gat, id_52gat, id_375gat);
and ( id_708gat, id_52gat, id_392gat);
and ( id_711gat, id_52gat, id_409gat);
and ( id_714gat, id_52gat, id_426gat);
and ( id_717gat, id_52gat, id_443gat);
and ( id_720gat, id_52gat, id_460gat);
and ( id_723gat, id_52gat, id_477gat);
and ( id_726gat, id_52gat, id_494gat);
and ( id_729gat, id_52gat, id_511gat);
and ( id_732gat, id_52gat, id_528gat);
and ( id_735gat, id_69gat, id_273gat);
and ( id_738gat, id_69gat, id_290gat);
and ( id_741gat, id_69gat, id_307gat);
and ( id_744gat, id_69gat, id_324gat);
and ( id_747gat, id_69gat, id_341gat);
and ( id_750gat, id_69gat, id_358gat);
and ( id_753gat, id_69gat, id_375gat);
and ( id_756gat, id_69gat, id_392gat);
and ( id_759gat, id_69gat, id_409gat);
and ( id_762gat, id_69gat, id_426gat);
and ( id_765gat, id_69gat, id_443gat);
and ( id_768gat, id_69gat, id_460gat);
and ( id_771gat, id_69gat, id_477gat);
and ( id_774gat, id_69gat, id_494gat);
and ( id_777gat, id_69gat, id_511gat);
and ( id_780gat, id_69gat, id_528gat);
and ( id_783gat, id_86gat, id_273gat);
and ( id_786gat, id_86gat, id_290gat);
and ( id_789gat, id_86gat, id_307gat);
and ( id_792gat, id_86gat, id_324gat);
and ( id_795gat, id_86gat, id_341gat);
and ( id_798gat, id_86gat, id_358gat);
and ( id_801gat, id_86gat, id_375gat);
and ( id_804gat, id_86gat, id_392gat);
and ( id_807gat, id_86gat, id_409gat);
and ( id_810gat, id_86gat, id_426gat);
and ( id_813gat, id_86gat, id_443gat);
and ( id_816gat, id_86gat, id_460gat);
and ( id_819gat, id_86gat, id_477gat);
and ( id_822gat, id_86gat, id_494gat);
and ( id_825gat, id_86gat, id_511gat);
and ( id_828gat, id_86gat, id_528gat);
and ( id_831gat, id_103gat, id_273gat);
and ( id_834gat, id_103gat, id_290gat);
and ( id_837gat, id_103gat, id_307gat);
and ( id_840gat, id_103gat, id_324gat);
and ( id_843gat, id_103gat, id_341gat);
and ( id_846gat, id_103gat, id_358gat);
and ( id_849gat, id_103gat, id_375gat);
and ( id_852gat, id_103gat, id_392gat);
and ( id_855gat, id_103gat, id_409gat);
and ( id_858gat, id_103gat, id_426gat);
and ( id_861gat, id_103gat, id_443gat);
and ( id_864gat, id_103gat, id_460gat);
and ( id_867gat, id_103gat, id_477gat);
and ( id_870gat, id_103gat, id_494gat);
and ( id_873gat, id_103gat, id_511gat);
and ( id_876gat, id_103gat, id_528gat);
and ( id_879gat, id_120gat, id_273gat);
and ( id_882gat, id_120gat, id_290gat);
and ( id_885gat, id_120gat, id_307gat);
and ( id_888gat, id_120gat, id_324gat);
and ( id_891gat, id_120gat, id_341gat);
and ( id_894gat, id_120gat, id_358gat);
and ( id_897gat, id_120gat, id_375gat);
and ( id_900gat, id_120gat, id_392gat);
and ( id_903gat, id_120gat, id_409gat);
and ( id_906gat, id_120gat, id_426gat);
and ( id_909gat, id_120gat, id_443gat);
and ( id_912gat, id_120gat, id_460gat);
and ( id_915gat, id_120gat, id_477gat);
and ( id_918gat, id_120gat, id_494gat);
and ( id_921gat, id_120gat, id_511gat);
and ( id_924gat, id_120gat, id_528gat);
and ( id_927gat, id_137gat, id_273gat);
and ( id_930gat, id_137gat, id_290gat);
and ( id_933gat, id_137gat, id_307gat);
and ( id_936gat, id_137gat, id_324gat);
and ( id_939gat, id_137gat, id_341gat);
and ( id_942gat, id_137gat, id_358gat);
and ( id_945gat, id_137gat, id_375gat);
and ( id_948gat, id_137gat, id_392gat);
and ( id_951gat, id_137gat, id_409gat);
and ( id_954gat, id_137gat, id_426gat);
and ( id_957gat, id_137gat, id_443gat);
and ( id_960gat, id_137gat, id_460gat);
and ( id_963gat, id_137gat, id_477gat);
and ( id_966gat, id_137gat, id_494gat);
and ( id_969gat, id_137gat, id_511gat);
and ( id_972gat, id_137gat, id_528gat);
and ( id_975gat, id_154gat, id_273gat);
and ( id_978gat, id_154gat, id_290gat);
and ( id_981gat, id_154gat, id_307gat);
and ( id_984gat, id_154gat, id_324gat);
and ( id_987gat, id_154gat, id_341gat);
and ( id_990gat, id_154gat, id_358gat);
and ( id_993gat, id_154gat, id_375gat);
and ( id_996gat, id_154gat, id_392gat);
and ( id_999gat, id_154gat, id_409gat);
and ( id_1002gat, id_154gat, id_426gat);
and ( id_1005gat, id_154gat, id_443gat);
and ( id_1008gat, id_154gat, id_460gat);
and ( id_1011gat, id_154gat, id_477gat);
and ( id_1014gat, id_154gat, id_494gat);
and ( id_1017gat, id_154gat, id_511gat);
and ( id_1020gat, id_154gat, id_528gat);
and ( id_1023gat, id_171gat, id_273gat);
and ( id_1026gat, id_171gat, id_290gat);
and ( id_1029gat, id_171gat, id_307gat);
and ( id_1032gat, id_171gat, id_324gat);
and ( id_1035gat, id_171gat, id_341gat);
and ( id_1038gat, id_171gat, id_358gat);
and ( id_1041gat, id_171gat, id_375gat);
and ( id_1044gat, id_171gat, id_392gat);
and ( id_1047gat, id_171gat, id_409gat);
and ( id_1050gat, id_171gat, id_426gat);
and ( id_1053gat, id_171gat, id_443gat);
and ( id_1056gat, id_171gat, id_460gat);
and ( id_1059gat, id_171gat, id_477gat);
and ( id_1062gat, id_171gat, id_494gat);
and ( id_1065gat, id_171gat, id_511gat);
and ( id_1068gat, id_171gat, id_528gat);
and ( id_1071gat, id_188gat, id_273gat);
and ( id_1074gat, id_188gat, id_290gat);
and ( id_1077gat, id_188gat, id_307gat);
and ( id_1080gat, id_188gat, id_324gat);
and ( id_1083gat, id_188gat, id_341gat);
and ( id_1086gat, id_188gat, id_358gat);
and ( id_1089gat, id_188gat, id_375gat);
and ( id_1092gat, id_188gat, id_392gat);
and ( id_1095gat, id_188gat, id_409gat);
and ( id_1098gat, id_188gat, id_426gat);
and ( id_1101gat, id_188gat, id_443gat);
and ( id_1104gat, id_188gat, id_460gat);
and ( id_1107gat, id_188gat, id_477gat);
and ( id_1110gat, id_188gat, id_494gat);
and ( id_1113gat, id_188gat, id_511gat);
and ( id_1116gat, id_188gat, id_528gat);
and ( id_1119gat, id_205gat, id_273gat);
and ( id_1122gat, id_205gat, id_290gat);
and ( id_1125gat, id_205gat, id_307gat);
and ( id_1128gat, id_205gat, id_324gat);
and ( id_1131gat, id_205gat, id_341gat);
and ( id_1134gat, id_205gat, id_358gat);
and ( id_1137gat, id_205gat, id_375gat);
and ( id_1140gat, id_205gat, id_392gat);
and ( id_1143gat, id_205gat, id_409gat);
and ( id_1146gat, id_205gat, id_426gat);
and ( id_1149gat, id_205gat, id_443gat);
and ( id_1152gat, id_205gat, id_460gat);
and ( id_1155gat, id_205gat, id_477gat);
and ( id_1158gat, id_205gat, id_494gat);
and ( id_1161gat, id_205gat, id_511gat);
and ( id_1164gat, id_205gat, id_528gat);
and ( id_1167gat, id_222gat, id_273gat);
and ( id_1170gat, id_222gat, id_290gat);
and ( id_1173gat, id_222gat, id_307gat);
and ( id_1176gat, id_222gat, id_324gat);
and ( id_1179gat, id_222gat, id_341gat);
and ( id_1182gat, id_222gat, id_358gat);
and ( id_1185gat, id_222gat, id_375gat);
and ( id_1188gat, id_222gat, id_392gat);
and ( id_1191gat, id_222gat, id_409gat);
and ( id_1194gat, id_222gat, id_426gat);
and ( id_1197gat, id_222gat, id_443gat);
and ( id_1200gat, id_222gat, id_460gat);
and ( id_1203gat, id_222gat, id_477gat);
and ( id_1206gat, id_222gat, id_494gat);
and ( id_1209gat, id_222gat, id_511gat);
and ( id_1212gat, id_222gat, id_528gat);
and ( id_1215gat, id_239gat, id_273gat);
and ( id_1218gat, id_239gat, id_290gat);
and ( id_1221gat, id_239gat, id_307gat);
and ( id_1224gat, id_239gat, id_324gat);
and ( id_1227gat, id_239gat, id_341gat);
and ( id_1230gat, id_239gat, id_358gat);
and ( id_1233gat, id_239gat, id_375gat);
and ( id_1236gat, id_239gat, id_392gat);
and ( id_1239gat, id_239gat, id_409gat);
and ( id_1242gat, id_239gat, id_426gat);
and ( id_1245gat, id_239gat, id_443gat);
and ( id_1248gat, id_239gat, id_460gat);
and ( id_1251gat, id_239gat, id_477gat);
and ( id_1254gat, id_239gat, id_494gat);
and ( id_1257gat, id_239gat, id_511gat);
and ( id_1260gat, id_239gat, id_528gat);
and ( id_1263gat, id_256gat, id_273gat);
and ( id_1266gat, id_256gat, id_290gat);
and ( id_1269gat, id_256gat, id_307gat);
and ( id_1272gat, id_256gat, id_324gat);
and ( id_1275gat, id_256gat, id_341gat);
and ( id_1278gat, id_256gat, id_358gat);
and ( id_1281gat, id_256gat, id_375gat);
and ( id_1284gat, id_256gat, id_392gat);
and ( id_1287gat, id_256gat, id_409gat);
and ( id_1290gat, id_256gat, id_426gat);
and ( id_1293gat, id_256gat, id_443gat);
and ( id_1296gat, id_256gat, id_460gat);
and ( id_1299gat, id_256gat, id_477gat);
and ( id_1302gat, id_256gat, id_494gat);
and ( id_1305gat, id_256gat, id_511gat);
and ( id_1308gat, id_256gat, id_528gat);
not ( id_1311gat, id_591gat);
not ( id_1315gat, id_639gat);
not ( id_1319gat, id_687gat);
not ( id_1323gat, id_735gat);
not ( id_1327gat, id_783gat);
not ( id_1331gat, id_831gat);
not ( id_1335gat, id_879gat);
not ( id_1339gat, id_927gat);
not ( id_1343gat, id_975gat);
not ( id_1347gat, id_1023gat);
not ( id_1351gat, id_1071gat);
not ( id_1355gat, id_1119gat);
not ( id_1359gat, id_1167gat);
not ( id_1363gat, id_1215gat);
not ( id_1367gat, id_1263gat);
not ( id_1372gat, id_1311gat);
not ( id_1374gat, id_1315gat);
not ( id_1376gat, id_1319gat);
not ( id_1378gat, id_1323gat);
not ( id_1380gat, id_1327gat);
not ( id_1382gat, id_1331gat);
not ( id_1384gat, id_1335gat);
not ( id_1386gat, id_1339gat);
not ( id_1388gat, id_1343gat);
not ( id_1390gat, id_1347gat);
not ( id_1392gat, id_1351gat);
not ( id_1394gat, id_1355gat);
not ( id_1396gat, id_1359gat);
not ( id_1398gat, id_1363gat);
not ( id_1400gat, id_1367gat);
not ( id_1401gat, id_1372gat);
not ( id_1404gat, id_1374gat);
not ( id_1407gat, id_1376gat);
not ( id_1410gat, id_1378gat);
not ( id_1413gat, id_1380gat);
not ( id_1416gat, id_1382gat);
not ( id_1419gat, id_1384gat);
not ( id_1422gat, id_1386gat);
not ( id_1425gat, id_1388gat);
not ( id_1428gat, id_1390gat);
not ( id_1431gat, id_1392gat);
not ( id_1434gat, id_1394gat);
not ( id_1437gat, id_1396gat);
not ( id_1440gat, id_1398gat);
not ( id_1443gat, id_1400gat);
nor ( id_1446gat, id_1401gat, id_546gat);
nor ( id_1450gat, id_1404gat, id_594gat);
nor ( id_1454gat, id_1407gat, id_642gat);
nor ( id_1458gat, id_1410gat, id_690gat);
nor ( id_1462gat, id_1413gat, id_738gat);
nor ( id_1466gat, id_1416gat, id_786gat);
nor ( id_1470gat, id_1419gat, id_834gat);
nor ( id_1474gat, id_1422gat, id_882gat);
nor ( id_1478gat, id_1425gat, id_930gat);
nor ( id_1482gat, id_1428gat, id_978gat);
nor ( id_1486gat, id_1431gat, id_1026gat);
nor ( id_1490gat, id_1434gat, id_1074gat);
nor ( id_1494gat, id_1437gat, id_1122gat);
nor ( id_1498gat, id_1440gat, id_1170gat);
nor ( id_1502gat, id_1443gat, id_1218gat);
nor ( id_1506gat, id_1401gat, id_1446gat);
nor ( id_1507gat, id_1446gat, id_546gat);
nor ( id_1508gat, id_1311gat, id_1446gat);
nor ( id_1511gat, id_1404gat, id_1450gat);
nor ( id_1512gat, id_1450gat, id_594gat);
nor ( id_1513gat, id_1315gat, id_1450gat);
nor ( id_1516gat, id_1407gat, id_1454gat);
nor ( id_1517gat, id_1454gat, id_642gat);
nor ( id_1518gat, id_1319gat, id_1454gat);
nor ( id_1521gat, id_1410gat, id_1458gat);
nor ( id_1522gat, id_1458gat, id_690gat);
nor ( id_1523gat, id_1323gat, id_1458gat);
nor ( id_1526gat, id_1413gat, id_1462gat);
nor ( id_1527gat, id_1462gat, id_738gat);
nor ( id_1528gat, id_1327gat, id_1462gat);
nor ( id_1531gat, id_1416gat, id_1466gat);
nor ( id_1532gat, id_1466gat, id_786gat);
nor ( id_1533gat, id_1331gat, id_1466gat);
nor ( id_1536gat, id_1419gat, id_1470gat);
nor ( id_1537gat, id_1470gat, id_834gat);
nor ( id_1538gat, id_1335gat, id_1470gat);
nor ( id_1541gat, id_1422gat, id_1474gat);
nor ( id_1542gat, id_1474gat, id_882gat);
nor ( id_1543gat, id_1339gat, id_1474gat);
nor ( id_1546gat, id_1425gat, id_1478gat);
nor ( id_1547gat, id_1478gat, id_930gat);
nor ( id_1548gat, id_1343gat, id_1478gat);
nor ( id_1551gat, id_1428gat, id_1482gat);
nor ( id_1552gat, id_1482gat, id_978gat);
nor ( id_1553gat, id_1347gat, id_1482gat);
nor ( id_1556gat, id_1431gat, id_1486gat);
nor ( id_1557gat, id_1486gat, id_1026gat);
nor ( id_1558gat, id_1351gat, id_1486gat);
nor ( id_1561gat, id_1434gat, id_1490gat);
nor ( id_1562gat, id_1490gat, id_1074gat);
nor ( id_1563gat, id_1355gat, id_1490gat);
nor ( id_1566gat, id_1437gat, id_1494gat);
nor ( id_1567gat, id_1494gat, id_1122gat);
nor ( id_1568gat, id_1359gat, id_1494gat);
nor ( id_1571gat, id_1440gat, id_1498gat);
nor ( id_1572gat, id_1498gat, id_1170gat);
nor ( id_1573gat, id_1363gat, id_1498gat);
nor ( id_1576gat, id_1443gat, id_1502gat);
nor ( id_1577gat, id_1502gat, id_1218gat);
nor ( id_1578gat, id_1367gat, id_1502gat);
nor ( id_1581gat, id_1506gat, id_1507gat);
nor ( id_1582gat, id_1511gat, id_1512gat);
nor ( id_1585gat, id_1516gat, id_1517gat);
nor ( id_1588gat, id_1521gat, id_1522gat);
nor ( id_1591gat, id_1526gat, id_1527gat);
nor ( id_1594gat, id_1531gat, id_1532gat);
nor ( id_1597gat, id_1536gat, id_1537gat);
nor ( id_1600gat, id_1541gat, id_1542gat);
nor ( id_1603gat, id_1546gat, id_1547gat);
nor ( id_1606gat, id_1551gat, id_1552gat);
nor ( id_1609gat, id_1556gat, id_1557gat);
nor ( id_1612gat, id_1561gat, id_1562gat);
nor ( id_1615gat, id_1566gat, id_1567gat);
nor ( id_1618gat, id_1571gat, id_1572gat);
nor ( id_1621gat, id_1576gat, id_1577gat);
not ( id_1624gat, id_1266gat);
nor ( id_1628gat, id_1582gat, id_1508gat);
nor ( id_1632gat, id_1585gat, id_1513gat);
nor ( id_1636gat, id_1588gat, id_1518gat);
nor ( id_1640gat, id_1591gat, id_1523gat);
nor ( id_1644gat, id_1594gat, id_1528gat);
nor ( id_1648gat, id_1597gat, id_1533gat);
nor ( id_1652gat, id_1600gat, id_1538gat);
nor ( id_1656gat, id_1603gat, id_1543gat);
nor ( id_1660gat, id_1606gat, id_1548gat);
nor ( id_1664gat, id_1609gat, id_1553gat);
nor ( id_1668gat, id_1612gat, id_1558gat);
nor ( id_1672gat, id_1615gat, id_1563gat);
nor ( id_1676gat, id_1618gat, id_1568gat);
nor ( id_1680gat, id_1621gat, id_1573gat);
nor ( id_1685gat, id_1624gat, id_1578gat);
nor ( id_1686gat, id_1582gat, id_1628gat);
nor ( id_1687gat, id_1628gat, id_1508gat);
nor ( id_1688gat, id_1585gat, id_1632gat);
nor ( id_1689gat, id_1632gat, id_1513gat);
nor ( id_1690gat, id_1588gat, id_1636gat);
nor ( id_1691gat, id_1636gat, id_1518gat);
nor ( id_1692gat, id_1591gat, id_1640gat);
nor ( id_1693gat, id_1640gat, id_1523gat);
nor ( id_1694gat, id_1594gat, id_1644gat);
nor ( id_1695gat, id_1644gat, id_1528gat);
nor ( id_1696gat, id_1597gat, id_1648gat);
nor ( id_1697gat, id_1648gat, id_1533gat);
nor ( id_1698gat, id_1600gat, id_1652gat);
nor ( id_1699gat, id_1652gat, id_1538gat);
nor ( id_1700gat, id_1603gat, id_1656gat);
nor ( id_1701gat, id_1656gat, id_1543gat);
nor ( id_1702gat, id_1606gat, id_1660gat);
nor ( id_1703gat, id_1660gat, id_1548gat);
nor ( id_1704gat, id_1609gat, id_1664gat);
nor ( id_1705gat, id_1664gat, id_1553gat);
nor ( id_1706gat, id_1612gat, id_1668gat);
nor ( id_1707gat, id_1668gat, id_1558gat);
nor ( id_1708gat, id_1615gat, id_1672gat);
nor ( id_1709gat, id_1672gat, id_1563gat);
nor ( id_1710gat, id_1618gat, id_1676gat);
nor ( id_1711gat, id_1676gat, id_1568gat);
nor ( id_1712gat, id_1621gat, id_1680gat);
nor ( id_1713gat, id_1680gat, id_1573gat);
not ( id_1714gat, id_1685gat);
nor ( id_1717gat, id_1686gat, id_1687gat);
nor ( id_1720gat, id_1688gat, id_1689gat);
nor ( id_1723gat, id_1690gat, id_1691gat);
nor ( id_1726gat, id_1692gat, id_1693gat);
nor ( id_1729gat, id_1694gat, id_1695gat);
nor ( id_1732gat, id_1696gat, id_1697gat);
nor ( id_1735gat, id_1698gat, id_1699gat);
nor ( id_1738gat, id_1700gat, id_1701gat);
nor ( id_1741gat, id_1702gat, id_1703gat);
nor ( id_1744gat, id_1704gat, id_1705gat);
nor ( id_1747gat, id_1706gat, id_1707gat);
nor ( id_1750gat, id_1708gat, id_1709gat);
nor ( id_1753gat, id_1710gat, id_1711gat);
nor ( id_1756gat, id_1712gat, id_1713gat);
nor ( id_1759gat, id_1714gat, id_1221gat);
nor ( id_1763gat, id_1717gat, id_549gat);
nor ( id_1767gat, id_1720gat, id_597gat);
nor ( id_1771gat, id_1723gat, id_645gat);
nor ( id_1775gat, id_1726gat, id_693gat);
nor ( id_1779gat, id_1729gat, id_741gat);
nor ( id_1783gat, id_1732gat, id_789gat);
nor ( id_1787gat, id_1735gat, id_837gat);
nor ( id_1791gat, id_1738gat, id_885gat);
nor ( id_1795gat, id_1741gat, id_933gat);
nor ( id_1799gat, id_1744gat, id_981gat);
nor ( id_1803gat, id_1747gat, id_1029gat);
nor ( id_1807gat, id_1750gat, id_1077gat);
nor ( id_1811gat, id_1753gat, id_1125gat);
nor ( id_1815gat, id_1756gat, id_1173gat);
nor ( id_1819gat, id_1714gat, id_1759gat);
nor ( id_1820gat, id_1759gat, id_1221gat);
nor ( id_1821gat, id_1624gat, id_1759gat);
nor ( id_1824gat, id_1717gat, id_1763gat);
nor ( id_1825gat, id_1763gat, id_549gat);
nor ( id_1826gat, id_1628gat, id_1763gat);
nor ( id_1829gat, id_1720gat, id_1767gat);
nor ( id_1830gat, id_1767gat, id_597gat);
nor ( id_1831gat, id_1632gat, id_1767gat);
nor ( id_1834gat, id_1723gat, id_1771gat);
nor ( id_1835gat, id_1771gat, id_645gat);
nor ( id_1836gat, id_1636gat, id_1771gat);
nor ( id_1839gat, id_1726gat, id_1775gat);
nor ( id_1840gat, id_1775gat, id_693gat);
nor ( id_1841gat, id_1640gat, id_1775gat);
nor ( id_1844gat, id_1729gat, id_1779gat);
nor ( id_1845gat, id_1779gat, id_741gat);
nor ( id_1846gat, id_1644gat, id_1779gat);
nor ( id_1849gat, id_1732gat, id_1783gat);
nor ( id_1850gat, id_1783gat, id_789gat);
nor ( id_1851gat, id_1648gat, id_1783gat);
nor ( id_1854gat, id_1735gat, id_1787gat);
nor ( id_1855gat, id_1787gat, id_837gat);
nor ( id_1856gat, id_1652gat, id_1787gat);
nor ( id_1859gat, id_1738gat, id_1791gat);
nor ( id_1860gat, id_1791gat, id_885gat);
nor ( id_1861gat, id_1656gat, id_1791gat);
nor ( id_1864gat, id_1741gat, id_1795gat);
nor ( id_1865gat, id_1795gat, id_933gat);
nor ( id_1866gat, id_1660gat, id_1795gat);
nor ( id_1869gat, id_1744gat, id_1799gat);
nor ( id_1870gat, id_1799gat, id_981gat);
nor ( id_1871gat, id_1664gat, id_1799gat);
nor ( id_1874gat, id_1747gat, id_1803gat);
nor ( id_1875gat, id_1803gat, id_1029gat);
nor ( id_1876gat, id_1668gat, id_1803gat);
nor ( id_1879gat, id_1750gat, id_1807gat);
nor ( id_1880gat, id_1807gat, id_1077gat);
nor ( id_1881gat, id_1672gat, id_1807gat);
nor ( id_1884gat, id_1753gat, id_1811gat);
nor ( id_1885gat, id_1811gat, id_1125gat);
nor ( id_1886gat, id_1676gat, id_1811gat);
nor ( id_1889gat, id_1756gat, id_1815gat);
nor ( id_1890gat, id_1815gat, id_1173gat);
nor ( id_1891gat, id_1680gat, id_1815gat);
nor ( id_1894gat, id_1819gat, id_1820gat);
nor ( id_1897gat, id_1269gat, id_1821gat);
nor ( id_1901gat, id_1824gat, id_1825gat);
nor ( id_1902gat, id_1829gat, id_1830gat);
nor ( id_1905gat, id_1834gat, id_1835gat);
nor ( id_1908gat, id_1839gat, id_1840gat);
nor ( id_1911gat, id_1844gat, id_1845gat);
nor ( id_1914gat, id_1849gat, id_1850gat);
nor ( id_1917gat, id_1854gat, id_1855gat);
nor ( id_1920gat, id_1859gat, id_1860gat);
nor ( id_1923gat, id_1864gat, id_1865gat);
nor ( id_1926gat, id_1869gat, id_1870gat);
nor ( id_1929gat, id_1874gat, id_1875gat);
nor ( id_1932gat, id_1879gat, id_1880gat);
nor ( id_1935gat, id_1884gat, id_1885gat);
nor ( id_1938gat, id_1889gat, id_1890gat);
nor ( id_1941gat, id_1894gat, id_1891gat);
nor ( id_1945gat, id_1269gat, id_1897gat);
nor ( id_1946gat, id_1897gat, id_1821gat);
nor ( id_1947gat, id_1902gat, id_1826gat);
nor ( id_1951gat, id_1905gat, id_1831gat);
nor ( id_1955gat, id_1908gat, id_1836gat);
nor ( id_1959gat, id_1911gat, id_1841gat);
nor ( id_1963gat, id_1914gat, id_1846gat);
nor ( id_1967gat, id_1917gat, id_1851gat);
nor ( id_1971gat, id_1920gat, id_1856gat);
nor ( id_1975gat, id_1923gat, id_1861gat);
nor ( id_1979gat, id_1926gat, id_1866gat);
nor ( id_1983gat, id_1929gat, id_1871gat);
nor ( id_1987gat, id_1932gat, id_1876gat);
nor ( id_1991gat, id_1935gat, id_1881gat);
nor ( id_1995gat, id_1938gat, id_1886gat);
nor ( id_1999gat, id_1894gat, id_1941gat);
nor ( id_2000gat, id_1941gat, id_1891gat);
nor ( id_2001gat, id_1945gat, id_1946gat);
nor ( id_2004gat, id_1902gat, id_1947gat);
nor ( id_2005gat, id_1947gat, id_1826gat);
nor ( id_2006gat, id_1905gat, id_1951gat);
nor ( id_2007gat, id_1951gat, id_1831gat);
nor ( id_2008gat, id_1908gat, id_1955gat);
nor ( id_2009gat, id_1955gat, id_1836gat);
nor ( id_2010gat, id_1911gat, id_1959gat);
nor ( id_2011gat, id_1959gat, id_1841gat);
nor ( id_2012gat, id_1914gat, id_1963gat);
nor ( id_2013gat, id_1963gat, id_1846gat);
nor ( id_2014gat, id_1917gat, id_1967gat);
nor ( id_2015gat, id_1967gat, id_1851gat);
nor ( id_2016gat, id_1920gat, id_1971gat);
nor ( id_2017gat, id_1971gat, id_1856gat);
nor ( id_2018gat, id_1923gat, id_1975gat);
nor ( id_2019gat, id_1975gat, id_1861gat);
nor ( id_2020gat, id_1926gat, id_1979gat);
nor ( id_2021gat, id_1979gat, id_1866gat);
nor ( id_2022gat, id_1929gat, id_1983gat);
nor ( id_2023gat, id_1983gat, id_1871gat);
nor ( id_2024gat, id_1932gat, id_1987gat);
nor ( id_2025gat, id_1987gat, id_1876gat);
nor ( id_2026gat, id_1935gat, id_1991gat);
nor ( id_2027gat, id_1991gat, id_1881gat);
nor ( id_2028gat, id_1938gat, id_1995gat);
nor ( id_2029gat, id_1995gat, id_1886gat);
nor ( id_2030gat, id_1999gat, id_2000gat);
nor ( id_2033gat, id_2001gat, id_1224gat);
nor ( id_2037gat, id_2004gat, id_2005gat);
nor ( id_2040gat, id_2006gat, id_2007gat);
nor ( id_2043gat, id_2008gat, id_2009gat);
nor ( id_2046gat, id_2010gat, id_2011gat);
nor ( id_2049gat, id_2012gat, id_2013gat);
nor ( id_2052gat, id_2014gat, id_2015gat);
nor ( id_2055gat, id_2016gat, id_2017gat);
nor ( id_2058gat, id_2018gat, id_2019gat);
nor ( id_2061gat, id_2020gat, id_2021gat);
nor ( id_2064gat, id_2022gat, id_2023gat);
nor ( id_2067gat, id_2024gat, id_2025gat);
nor ( id_2070gat, id_2026gat, id_2027gat);
nor ( id_2073gat, id_2028gat, id_2029gat);
nor ( id_2076gat, id_2030gat, id_1176gat);
nor ( id_2080gat, id_2001gat, id_2033gat);
nor ( id_2081gat, id_2033gat, id_1224gat);
nor ( id_2082gat, id_1897gat, id_2033gat);
nor ( id_2085gat, id_2037gat, id_552gat);
nor ( id_2089gat, id_2040gat, id_600gat);
nor ( id_2093gat, id_2043gat, id_648gat);
nor ( id_2097gat, id_2046gat, id_696gat);
nor ( id_2101gat, id_2049gat, id_744gat);
nor ( id_2105gat, id_2052gat, id_792gat);
nor ( id_2109gat, id_2055gat, id_840gat);
nor ( id_2113gat, id_2058gat, id_888gat);
nor ( id_2117gat, id_2061gat, id_936gat);
nor ( id_2121gat, id_2064gat, id_984gat);
nor ( id_2125gat, id_2067gat, id_1032gat);
nor ( id_2129gat, id_2070gat, id_1080gat);
nor ( id_2133gat, id_2073gat, id_1128gat);
nor ( id_2137gat, id_2030gat, id_2076gat);
nor ( id_2138gat, id_2076gat, id_1176gat);
nor ( id_2139gat, id_1941gat, id_2076gat);
nor ( id_2142gat, id_2080gat, id_2081gat);
nor ( id_2145gat, id_1272gat, id_2082gat);
nor ( id_2149gat, id_2037gat, id_2085gat);
nor ( id_2150gat, id_2085gat, id_552gat);
nor ( id_2151gat, id_1947gat, id_2085gat);
nor ( id_2154gat, id_2040gat, id_2089gat);
nor ( id_2155gat, id_2089gat, id_600gat);
nor ( id_2156gat, id_1951gat, id_2089gat);
nor ( id_2159gat, id_2043gat, id_2093gat);
nor ( id_2160gat, id_2093gat, id_648gat);
nor ( id_2161gat, id_1955gat, id_2093gat);
nor ( id_2164gat, id_2046gat, id_2097gat);
nor ( id_2165gat, id_2097gat, id_696gat);
nor ( id_2166gat, id_1959gat, id_2097gat);
nor ( id_2169gat, id_2049gat, id_2101gat);
nor ( id_2170gat, id_2101gat, id_744gat);
nor ( id_2171gat, id_1963gat, id_2101gat);
nor ( id_2174gat, id_2052gat, id_2105gat);
nor ( id_2175gat, id_2105gat, id_792gat);
nor ( id_2176gat, id_1967gat, id_2105gat);
nor ( id_2179gat, id_2055gat, id_2109gat);
nor ( id_2180gat, id_2109gat, id_840gat);
nor ( id_2181gat, id_1971gat, id_2109gat);
nor ( id_2184gat, id_2058gat, id_2113gat);
nor ( id_2185gat, id_2113gat, id_888gat);
nor ( id_2186gat, id_1975gat, id_2113gat);
nor ( id_2189gat, id_2061gat, id_2117gat);
nor ( id_2190gat, id_2117gat, id_936gat);
nor ( id_2191gat, id_1979gat, id_2117gat);
nor ( id_2194gat, id_2064gat, id_2121gat);
nor ( id_2195gat, id_2121gat, id_984gat);
nor ( id_2196gat, id_1983gat, id_2121gat);
nor ( id_2199gat, id_2067gat, id_2125gat);
nor ( id_2200gat, id_2125gat, id_1032gat);
nor ( id_2201gat, id_1987gat, id_2125gat);
nor ( id_2204gat, id_2070gat, id_2129gat);
nor ( id_2205gat, id_2129gat, id_1080gat);
nor ( id_2206gat, id_1991gat, id_2129gat);
nor ( id_2209gat, id_2073gat, id_2133gat);
nor ( id_2210gat, id_2133gat, id_1128gat);
nor ( id_2211gat, id_1995gat, id_2133gat);
nor ( id_2214gat, id_2137gat, id_2138gat);
nor ( id_2217gat, id_2142gat, id_2139gat);
nor ( id_2221gat, id_1272gat, id_2145gat);
nor ( id_2222gat, id_2145gat, id_2082gat);
nor ( id_2223gat, id_2149gat, id_2150gat);
nor ( id_2224gat, id_2154gat, id_2155gat);
nor ( id_2227gat, id_2159gat, id_2160gat);
nor ( id_2230gat, id_2164gat, id_2165gat);
nor ( id_2233gat, id_2169gat, id_2170gat);
nor ( id_2236gat, id_2174gat, id_2175gat);
nor ( id_2239gat, id_2179gat, id_2180gat);
nor ( id_2242gat, id_2184gat, id_2185gat);
nor ( id_2245gat, id_2189gat, id_2190gat);
nor ( id_2248gat, id_2194gat, id_2195gat);
nor ( id_2251gat, id_2199gat, id_2200gat);
nor ( id_2254gat, id_2204gat, id_2205gat);
nor ( id_2257gat, id_2209gat, id_2210gat);
nor ( id_2260gat, id_2214gat, id_2211gat);
nor ( id_2264gat, id_2142gat, id_2217gat);
nor ( id_2265gat, id_2217gat, id_2139gat);
nor ( id_2266gat, id_2221gat, id_2222gat);
nor ( id_2269gat, id_2224gat, id_2151gat);
nor ( id_2273gat, id_2227gat, id_2156gat);
nor ( id_2277gat, id_2230gat, id_2161gat);
nor ( id_2281gat, id_2233gat, id_2166gat);
nor ( id_2285gat, id_2236gat, id_2171gat);
nor ( id_2289gat, id_2239gat, id_2176gat);
nor ( id_2293gat, id_2242gat, id_2181gat);
nor ( id_2297gat, id_2245gat, id_2186gat);
nor ( id_2301gat, id_2248gat, id_2191gat);
nor ( id_2305gat, id_2251gat, id_2196gat);
nor ( id_2309gat, id_2254gat, id_2201gat);
nor ( id_2313gat, id_2257gat, id_2206gat);
nor ( id_2317gat, id_2214gat, id_2260gat);
nor ( id_2318gat, id_2260gat, id_2211gat);
nor ( id_2319gat, id_2264gat, id_2265gat);
nor ( id_2322gat, id_2266gat, id_1227gat);
nor ( id_2326gat, id_2224gat, id_2269gat);
nor ( id_2327gat, id_2269gat, id_2151gat);
nor ( id_2328gat, id_2227gat, id_2273gat);
nor ( id_2329gat, id_2273gat, id_2156gat);
nor ( id_2330gat, id_2230gat, id_2277gat);
nor ( id_2331gat, id_2277gat, id_2161gat);
nor ( id_2332gat, id_2233gat, id_2281gat);
nor ( id_2333gat, id_2281gat, id_2166gat);
nor ( id_2334gat, id_2236gat, id_2285gat);
nor ( id_2335gat, id_2285gat, id_2171gat);
nor ( id_2336gat, id_2239gat, id_2289gat);
nor ( id_2337gat, id_2289gat, id_2176gat);
nor ( id_2338gat, id_2242gat, id_2293gat);
nor ( id_2339gat, id_2293gat, id_2181gat);
nor ( id_2340gat, id_2245gat, id_2297gat);
nor ( id_2341gat, id_2297gat, id_2186gat);
nor ( id_2342gat, id_2248gat, id_2301gat);
nor ( id_2343gat, id_2301gat, id_2191gat);
nor ( id_2344gat, id_2251gat, id_2305gat);
nor ( id_2345gat, id_2305gat, id_2196gat);
nor ( id_2346gat, id_2254gat, id_2309gat);
nor ( id_2347gat, id_2309gat, id_2201gat);
nor ( id_2348gat, id_2257gat, id_2313gat);
nor ( id_2349gat, id_2313gat, id_2206gat);
nor ( id_2350gat, id_2317gat, id_2318gat);
nor ( id_2353gat, id_2319gat, id_1179gat);
nor ( id_2357gat, id_2266gat, id_2322gat);
nor ( id_2358gat, id_2322gat, id_1227gat);
nor ( id_2359gat, id_2145gat, id_2322gat);
nor ( id_2362gat, id_2326gat, id_2327gat);
nor ( id_2365gat, id_2328gat, id_2329gat);
nor ( id_2368gat, id_2330gat, id_2331gat);
nor ( id_2371gat, id_2332gat, id_2333gat);
nor ( id_2374gat, id_2334gat, id_2335gat);
nor ( id_2377gat, id_2336gat, id_2337gat);
nor ( id_2380gat, id_2338gat, id_2339gat);
nor ( id_2383gat, id_2340gat, id_2341gat);
nor ( id_2386gat, id_2342gat, id_2343gat);
nor ( id_2389gat, id_2344gat, id_2345gat);
nor ( id_2392gat, id_2346gat, id_2347gat);
nor ( id_2395gat, id_2348gat, id_2349gat);
nor ( id_2398gat, id_2350gat, id_1131gat);
nor ( id_2402gat, id_2319gat, id_2353gat);
nor ( id_2403gat, id_2353gat, id_1179gat);
nor ( id_2404gat, id_2217gat, id_2353gat);
nor ( id_2407gat, id_2357gat, id_2358gat);
nor ( id_2410gat, id_1275gat, id_2359gat);
nor ( id_2414gat, id_2362gat, id_555gat);
nor ( id_2418gat, id_2365gat, id_603gat);
nor ( id_2422gat, id_2368gat, id_651gat);
nor ( id_2426gat, id_2371gat, id_699gat);
nor ( id_2430gat, id_2374gat, id_747gat);
nor ( id_2434gat, id_2377gat, id_795gat);
nor ( id_2438gat, id_2380gat, id_843gat);
nor ( id_2442gat, id_2383gat, id_891gat);
nor ( id_2446gat, id_2386gat, id_939gat);
nor ( id_2450gat, id_2389gat, id_987gat);
nor ( id_2454gat, id_2392gat, id_1035gat);
nor ( id_2458gat, id_2395gat, id_1083gat);
nor ( id_2462gat, id_2350gat, id_2398gat);
nor ( id_2463gat, id_2398gat, id_1131gat);
nor ( id_2464gat, id_2260gat, id_2398gat);
nor ( id_2467gat, id_2402gat, id_2403gat);
nor ( id_2470gat, id_2407gat, id_2404gat);
nor ( id_2474gat, id_1275gat, id_2410gat);
nor ( id_2475gat, id_2410gat, id_2359gat);
nor ( id_2476gat, id_2362gat, id_2414gat);
nor ( id_2477gat, id_2414gat, id_555gat);
nor ( id_2478gat, id_2269gat, id_2414gat);
nor ( id_2481gat, id_2365gat, id_2418gat);
nor ( id_2482gat, id_2418gat, id_603gat);
nor ( id_2483gat, id_2273gat, id_2418gat);
nor ( id_2486gat, id_2368gat, id_2422gat);
nor ( id_2487gat, id_2422gat, id_651gat);
nor ( id_2488gat, id_2277gat, id_2422gat);
nor ( id_2491gat, id_2371gat, id_2426gat);
nor ( id_2492gat, id_2426gat, id_699gat);
nor ( id_2493gat, id_2281gat, id_2426gat);
nor ( id_2496gat, id_2374gat, id_2430gat);
nor ( id_2497gat, id_2430gat, id_747gat);
nor ( id_2498gat, id_2285gat, id_2430gat);
nor ( id_2501gat, id_2377gat, id_2434gat);
nor ( id_2502gat, id_2434gat, id_795gat);
nor ( id_2503gat, id_2289gat, id_2434gat);
nor ( id_2506gat, id_2380gat, id_2438gat);
nor ( id_2507gat, id_2438gat, id_843gat);
nor ( id_2508gat, id_2293gat, id_2438gat);
nor ( id_2511gat, id_2383gat, id_2442gat);
nor ( id_2512gat, id_2442gat, id_891gat);
nor ( id_2513gat, id_2297gat, id_2442gat);
nor ( id_2516gat, id_2386gat, id_2446gat);
nor ( id_2517gat, id_2446gat, id_939gat);
nor ( id_2518gat, id_2301gat, id_2446gat);
nor ( id_2521gat, id_2389gat, id_2450gat);
nor ( id_2522gat, id_2450gat, id_987gat);
nor ( id_2523gat, id_2305gat, id_2450gat);
nor ( id_2526gat, id_2392gat, id_2454gat);
nor ( id_2527gat, id_2454gat, id_1035gat);
nor ( id_2528gat, id_2309gat, id_2454gat);
nor ( id_2531gat, id_2395gat, id_2458gat);
nor ( id_2532gat, id_2458gat, id_1083gat);
nor ( id_2533gat, id_2313gat, id_2458gat);
nor ( id_2536gat, id_2462gat, id_2463gat);
nor ( id_2539gat, id_2467gat, id_2464gat);
nor ( id_2543gat, id_2407gat, id_2470gat);
nor ( id_2544gat, id_2470gat, id_2404gat);
nor ( id_2545gat, id_2474gat, id_2475gat);
nor ( id_2548gat, id_2476gat, id_2477gat);
nor ( id_2549gat, id_2481gat, id_2482gat);
nor ( id_2552gat, id_2486gat, id_2487gat);
nor ( id_2555gat, id_2491gat, id_2492gat);
nor ( id_2558gat, id_2496gat, id_2497gat);
nor ( id_2561gat, id_2501gat, id_2502gat);
nor ( id_2564gat, id_2506gat, id_2507gat);
nor ( id_2567gat, id_2511gat, id_2512gat);
nor ( id_2570gat, id_2516gat, id_2517gat);
nor ( id_2573gat, id_2521gat, id_2522gat);
nor ( id_2576gat, id_2526gat, id_2527gat);
nor ( id_2579gat, id_2531gat, id_2532gat);
nor ( id_2582gat, id_2536gat, id_2533gat);
nor ( id_2586gat, id_2467gat, id_2539gat);
nor ( id_2587gat, id_2539gat, id_2464gat);
nor ( id_2588gat, id_2543gat, id_2544gat);
nor ( id_2591gat, id_2545gat, id_1230gat);
nor ( id_2595gat, id_2549gat, id_2478gat);
nor ( id_2599gat, id_2552gat, id_2483gat);
nor ( id_2603gat, id_2555gat, id_2488gat);
nor ( id_2607gat, id_2558gat, id_2493gat);
nor ( id_2611gat, id_2561gat, id_2498gat);
nor ( id_2615gat, id_2564gat, id_2503gat);
nor ( id_2619gat, id_2567gat, id_2508gat);
nor ( id_2623gat, id_2570gat, id_2513gat);
nor ( id_2627gat, id_2573gat, id_2518gat);
nor ( id_2631gat, id_2576gat, id_2523gat);
nor ( id_2635gat, id_2579gat, id_2528gat);
nor ( id_2639gat, id_2536gat, id_2582gat);
nor ( id_2640gat, id_2582gat, id_2533gat);
nor ( id_2641gat, id_2586gat, id_2587gat);
nor ( id_2644gat, id_2588gat, id_1182gat);
nor ( id_2648gat, id_2545gat, id_2591gat);
nor ( id_2649gat, id_2591gat, id_1230gat);
nor ( id_2650gat, id_2410gat, id_2591gat);
nor ( id_2653gat, id_2549gat, id_2595gat);
nor ( id_2654gat, id_2595gat, id_2478gat);
nor ( id_2655gat, id_2552gat, id_2599gat);
nor ( id_2656gat, id_2599gat, id_2483gat);
nor ( id_2657gat, id_2555gat, id_2603gat);
nor ( id_2658gat, id_2603gat, id_2488gat);
nor ( id_2659gat, id_2558gat, id_2607gat);
nor ( id_2660gat, id_2607gat, id_2493gat);
nor ( id_2661gat, id_2561gat, id_2611gat);
nor ( id_2662gat, id_2611gat, id_2498gat);
nor ( id_2663gat, id_2564gat, id_2615gat);
nor ( id_2664gat, id_2615gat, id_2503gat);
nor ( id_2665gat, id_2567gat, id_2619gat);
nor ( id_2666gat, id_2619gat, id_2508gat);
nor ( id_2667gat, id_2570gat, id_2623gat);
nor ( id_2668gat, id_2623gat, id_2513gat);
nor ( id_2669gat, id_2573gat, id_2627gat);
nor ( id_2670gat, id_2627gat, id_2518gat);
nor ( id_2671gat, id_2576gat, id_2631gat);
nor ( id_2672gat, id_2631gat, id_2523gat);
nor ( id_2673gat, id_2579gat, id_2635gat);
nor ( id_2674gat, id_2635gat, id_2528gat);
nor ( id_2675gat, id_2639gat, id_2640gat);
nor ( id_2678gat, id_2641gat, id_1134gat);
nor ( id_2682gat, id_2588gat, id_2644gat);
nor ( id_2683gat, id_2644gat, id_1182gat);
nor ( id_2684gat, id_2470gat, id_2644gat);
nor ( id_2687gat, id_2648gat, id_2649gat);
nor ( id_2690gat, id_1278gat, id_2650gat);
nor ( id_2694gat, id_2653gat, id_2654gat);
nor ( id_2697gat, id_2655gat, id_2656gat);
nor ( id_2700gat, id_2657gat, id_2658gat);
nor ( id_2703gat, id_2659gat, id_2660gat);
nor ( id_2706gat, id_2661gat, id_2662gat);
nor ( id_2709gat, id_2663gat, id_2664gat);
nor ( id_2712gat, id_2665gat, id_2666gat);
nor ( id_2715gat, id_2667gat, id_2668gat);
nor ( id_2718gat, id_2669gat, id_2670gat);
nor ( id_2721gat, id_2671gat, id_2672gat);
nor ( id_2724gat, id_2673gat, id_2674gat);
nor ( id_2727gat, id_2675gat, id_1086gat);
nor ( id_2731gat, id_2641gat, id_2678gat);
nor ( id_2732gat, id_2678gat, id_1134gat);
nor ( id_2733gat, id_2539gat, id_2678gat);
nor ( id_2736gat, id_2682gat, id_2683gat);
nor ( id_2739gat, id_2687gat, id_2684gat);
nor ( id_2743gat, id_1278gat, id_2690gat);
nor ( id_2744gat, id_2690gat, id_2650gat);
nor ( id_2745gat, id_2694gat, id_558gat);
nor ( id_2749gat, id_2697gat, id_606gat);
nor ( id_2753gat, id_2700gat, id_654gat);
nor ( id_2757gat, id_2703gat, id_702gat);
nor ( id_2761gat, id_2706gat, id_750gat);
nor ( id_2765gat, id_2709gat, id_798gat);
nor ( id_2769gat, id_2712gat, id_846gat);
nor ( id_2773gat, id_2715gat, id_894gat);
nor ( id_2777gat, id_2718gat, id_942gat);
nor ( id_2781gat, id_2721gat, id_990gat);
nor ( id_2785gat, id_2724gat, id_1038gat);
nor ( id_2789gat, id_2675gat, id_2727gat);
nor ( id_2790gat, id_2727gat, id_1086gat);
nor ( id_2791gat, id_2582gat, id_2727gat);
nor ( id_2794gat, id_2731gat, id_2732gat);
nor ( id_2797gat, id_2736gat, id_2733gat);
nor ( id_2801gat, id_2687gat, id_2739gat);
nor ( id_2802gat, id_2739gat, id_2684gat);
nor ( id_2803gat, id_2743gat, id_2744gat);
nor ( id_2806gat, id_2694gat, id_2745gat);
nor ( id_2807gat, id_2745gat, id_558gat);
nor ( id_2808gat, id_2595gat, id_2745gat);
nor ( id_2811gat, id_2697gat, id_2749gat);
nor ( id_2812gat, id_2749gat, id_606gat);
nor ( id_2813gat, id_2599gat, id_2749gat);
nor ( id_2816gat, id_2700gat, id_2753gat);
nor ( id_2817gat, id_2753gat, id_654gat);
nor ( id_2818gat, id_2603gat, id_2753gat);
nor ( id_2821gat, id_2703gat, id_2757gat);
nor ( id_2822gat, id_2757gat, id_702gat);
nor ( id_2823gat, id_2607gat, id_2757gat);
nor ( id_2826gat, id_2706gat, id_2761gat);
nor ( id_2827gat, id_2761gat, id_750gat);
nor ( id_2828gat, id_2611gat, id_2761gat);
nor ( id_2831gat, id_2709gat, id_2765gat);
nor ( id_2832gat, id_2765gat, id_798gat);
nor ( id_2833gat, id_2615gat, id_2765gat);
nor ( id_2836gat, id_2712gat, id_2769gat);
nor ( id_2837gat, id_2769gat, id_846gat);
nor ( id_2838gat, id_2619gat, id_2769gat);
nor ( id_2841gat, id_2715gat, id_2773gat);
nor ( id_2842gat, id_2773gat, id_894gat);
nor ( id_2843gat, id_2623gat, id_2773gat);
nor ( id_2846gat, id_2718gat, id_2777gat);
nor ( id_2847gat, id_2777gat, id_942gat);
nor ( id_2848gat, id_2627gat, id_2777gat);
nor ( id_2851gat, id_2721gat, id_2781gat);
nor ( id_2852gat, id_2781gat, id_990gat);
nor ( id_2853gat, id_2631gat, id_2781gat);
nor ( id_2856gat, id_2724gat, id_2785gat);
nor ( id_2857gat, id_2785gat, id_1038gat);
nor ( id_2858gat, id_2635gat, id_2785gat);
nor ( id_2861gat, id_2789gat, id_2790gat);
nor ( id_2864gat, id_2794gat, id_2791gat);
nor ( id_2868gat, id_2736gat, id_2797gat);
nor ( id_2869gat, id_2797gat, id_2733gat);
nor ( id_2870gat, id_2801gat, id_2802gat);
nor ( id_2873gat, id_2803gat, id_1233gat);
nor ( id_2877gat, id_2806gat, id_2807gat);
nor ( id_2878gat, id_2811gat, id_2812gat);
nor ( id_2881gat, id_2816gat, id_2817gat);
nor ( id_2884gat, id_2821gat, id_2822gat);
nor ( id_2887gat, id_2826gat, id_2827gat);
nor ( id_2890gat, id_2831gat, id_2832gat);
nor ( id_2893gat, id_2836gat, id_2837gat);
nor ( id_2896gat, id_2841gat, id_2842gat);
nor ( id_2899gat, id_2846gat, id_2847gat);
nor ( id_2902gat, id_2851gat, id_2852gat);
nor ( id_2905gat, id_2856gat, id_2857gat);
nor ( id_2908gat, id_2861gat, id_2858gat);
nor ( id_2912gat, id_2794gat, id_2864gat);
nor ( id_2913gat, id_2864gat, id_2791gat);
nor ( id_2914gat, id_2868gat, id_2869gat);
nor ( id_2917gat, id_2870gat, id_1185gat);
nor ( id_2921gat, id_2803gat, id_2873gat);
nor ( id_2922gat, id_2873gat, id_1233gat);
nor ( id_2923gat, id_2690gat, id_2873gat);
nor ( id_2926gat, id_2878gat, id_2808gat);
nor ( id_2930gat, id_2881gat, id_2813gat);
nor ( id_2934gat, id_2884gat, id_2818gat);
nor ( id_2938gat, id_2887gat, id_2823gat);
nor ( id_2942gat, id_2890gat, id_2828gat);
nor ( id_2946gat, id_2893gat, id_2833gat);
nor ( id_2950gat, id_2896gat, id_2838gat);
nor ( id_2954gat, id_2899gat, id_2843gat);
nor ( id_2958gat, id_2902gat, id_2848gat);
nor ( id_2962gat, id_2905gat, id_2853gat);
nor ( id_2966gat, id_2861gat, id_2908gat);
nor ( id_2967gat, id_2908gat, id_2858gat);
nor ( id_2968gat, id_2912gat, id_2913gat);
nor ( id_2971gat, id_2914gat, id_1137gat);
nor ( id_2975gat, id_2870gat, id_2917gat);
nor ( id_2976gat, id_2917gat, id_1185gat);
nor ( id_2977gat, id_2739gat, id_2917gat);
nor ( id_2980gat, id_2921gat, id_2922gat);
nor ( id_2983gat, id_1281gat, id_2923gat);
nor ( id_2987gat, id_2878gat, id_2926gat);
nor ( id_2988gat, id_2926gat, id_2808gat);
nor ( id_2989gat, id_2881gat, id_2930gat);
nor ( id_2990gat, id_2930gat, id_2813gat);
nor ( id_2991gat, id_2884gat, id_2934gat);
nor ( id_2992gat, id_2934gat, id_2818gat);
nor ( id_2993gat, id_2887gat, id_2938gat);
nor ( id_2994gat, id_2938gat, id_2823gat);
nor ( id_2995gat, id_2890gat, id_2942gat);
nor ( id_2996gat, id_2942gat, id_2828gat);
nor ( id_2997gat, id_2893gat, id_2946gat);
nor ( id_2998gat, id_2946gat, id_2833gat);
nor ( id_2999gat, id_2896gat, id_2950gat);
nor ( id_3000gat, id_2950gat, id_2838gat);
nor ( id_3001gat, id_2899gat, id_2954gat);
nor ( id_3002gat, id_2954gat, id_2843gat);
nor ( id_3003gat, id_2902gat, id_2958gat);
nor ( id_3004gat, id_2958gat, id_2848gat);
nor ( id_3005gat, id_2905gat, id_2962gat);
nor ( id_3006gat, id_2962gat, id_2853gat);
nor ( id_3007gat, id_2966gat, id_2967gat);
nor ( id_3010gat, id_2968gat, id_1089gat);
nor ( id_3014gat, id_2914gat, id_2971gat);
nor ( id_3015gat, id_2971gat, id_1137gat);
nor ( id_3016gat, id_2797gat, id_2971gat);
nor ( id_3019gat, id_2975gat, id_2976gat);
nor ( id_3022gat, id_2980gat, id_2977gat);
nor ( id_3026gat, id_1281gat, id_2983gat);
nor ( id_3027gat, id_2983gat, id_2923gat);
nor ( id_3028gat, id_2987gat, id_2988gat);
nor ( id_3031gat, id_2989gat, id_2990gat);
nor ( id_3034gat, id_2991gat, id_2992gat);
nor ( id_3037gat, id_2993gat, id_2994gat);
nor ( id_3040gat, id_2995gat, id_2996gat);
nor ( id_3043gat, id_2997gat, id_2998gat);
nor ( id_3046gat, id_2999gat, id_3000gat);
nor ( id_3049gat, id_3001gat, id_3002gat);
nor ( id_3052gat, id_3003gat, id_3004gat);
nor ( id_3055gat, id_3005gat, id_3006gat);
nor ( id_3058gat, id_3007gat, id_1041gat);
nor ( id_3062gat, id_2968gat, id_3010gat);
nor ( id_3063gat, id_3010gat, id_1089gat);
nor ( id_3064gat, id_2864gat, id_3010gat);
nor ( id_3067gat, id_3014gat, id_3015gat);
nor ( id_3070gat, id_3019gat, id_3016gat);
nor ( id_3074gat, id_2980gat, id_3022gat);
nor ( id_3075gat, id_3022gat, id_2977gat);
nor ( id_3076gat, id_3026gat, id_3027gat);
nor ( id_3079gat, id_3028gat, id_561gat);
nor ( id_3083gat, id_3031gat, id_609gat);
nor ( id_3087gat, id_3034gat, id_657gat);
nor ( id_3091gat, id_3037gat, id_705gat);
nor ( id_3095gat, id_3040gat, id_753gat);
nor ( id_3099gat, id_3043gat, id_801gat);
nor ( id_3103gat, id_3046gat, id_849gat);
nor ( id_3107gat, id_3049gat, id_897gat);
nor ( id_3111gat, id_3052gat, id_945gat);
nor ( id_3115gat, id_3055gat, id_993gat);
nor ( id_3119gat, id_3007gat, id_3058gat);
nor ( id_3120gat, id_3058gat, id_1041gat);
nor ( id_3121gat, id_2908gat, id_3058gat);
nor ( id_3124gat, id_3062gat, id_3063gat);
nor ( id_3127gat, id_3067gat, id_3064gat);
nor ( id_3131gat, id_3019gat, id_3070gat);
nor ( id_3132gat, id_3070gat, id_3016gat);
nor ( id_3133gat, id_3074gat, id_3075gat);
nor ( id_3136gat, id_3076gat, id_1236gat);
nor ( id_3140gat, id_3028gat, id_3079gat);
nor ( id_3141gat, id_3079gat, id_561gat);
nor ( id_3142gat, id_2926gat, id_3079gat);
nor ( id_3145gat, id_3031gat, id_3083gat);
nor ( id_3146gat, id_3083gat, id_609gat);
nor ( id_3147gat, id_2930gat, id_3083gat);
nor ( id_3150gat, id_3034gat, id_3087gat);
nor ( id_3151gat, id_3087gat, id_657gat);
nor ( id_3152gat, id_2934gat, id_3087gat);
nor ( id_3155gat, id_3037gat, id_3091gat);
nor ( id_3156gat, id_3091gat, id_705gat);
nor ( id_3157gat, id_2938gat, id_3091gat);
nor ( id_3160gat, id_3040gat, id_3095gat);
nor ( id_3161gat, id_3095gat, id_753gat);
nor ( id_3162gat, id_2942gat, id_3095gat);
nor ( id_3165gat, id_3043gat, id_3099gat);
nor ( id_3166gat, id_3099gat, id_801gat);
nor ( id_3167gat, id_2946gat, id_3099gat);
nor ( id_3170gat, id_3046gat, id_3103gat);
nor ( id_3171gat, id_3103gat, id_849gat);
nor ( id_3172gat, id_2950gat, id_3103gat);
nor ( id_3175gat, id_3049gat, id_3107gat);
nor ( id_3176gat, id_3107gat, id_897gat);
nor ( id_3177gat, id_2954gat, id_3107gat);
nor ( id_3180gat, id_3052gat, id_3111gat);
nor ( id_3181gat, id_3111gat, id_945gat);
nor ( id_3182gat, id_2958gat, id_3111gat);
nor ( id_3185gat, id_3055gat, id_3115gat);
nor ( id_3186gat, id_3115gat, id_993gat);
nor ( id_3187gat, id_2962gat, id_3115gat);
nor ( id_3190gat, id_3119gat, id_3120gat);
nor ( id_3193gat, id_3124gat, id_3121gat);
nor ( id_3197gat, id_3067gat, id_3127gat);
nor ( id_3198gat, id_3127gat, id_3064gat);
nor ( id_3199gat, id_3131gat, id_3132gat);
nor ( id_3202gat, id_3133gat, id_1188gat);
nor ( id_3206gat, id_3076gat, id_3136gat);
nor ( id_3207gat, id_3136gat, id_1236gat);
nor ( id_3208gat, id_2983gat, id_3136gat);
nor ( id_3211gat, id_3140gat, id_3141gat);
nor ( id_3212gat, id_3145gat, id_3146gat);
nor ( id_3215gat, id_3150gat, id_3151gat);
nor ( id_3218gat, id_3155gat, id_3156gat);
nor ( id_3221gat, id_3160gat, id_3161gat);
nor ( id_3224gat, id_3165gat, id_3166gat);
nor ( id_3227gat, id_3170gat, id_3171gat);
nor ( id_3230gat, id_3175gat, id_3176gat);
nor ( id_3233gat, id_3180gat, id_3181gat);
nor ( id_3236gat, id_3185gat, id_3186gat);
nor ( id_3239gat, id_3190gat, id_3187gat);
nor ( id_3243gat, id_3124gat, id_3193gat);
nor ( id_3244gat, id_3193gat, id_3121gat);
nor ( id_3245gat, id_3197gat, id_3198gat);
nor ( id_3248gat, id_3199gat, id_1140gat);
nor ( id_3252gat, id_3133gat, id_3202gat);
nor ( id_3253gat, id_3202gat, id_1188gat);
nor ( id_3254gat, id_3022gat, id_3202gat);
nor ( id_3257gat, id_3206gat, id_3207gat);
nor ( id_3260gat, id_1284gat, id_3208gat);
nor ( id_3264gat, id_3212gat, id_3142gat);
nor ( id_3268gat, id_3215gat, id_3147gat);
nor ( id_3272gat, id_3218gat, id_3152gat);
nor ( id_3276gat, id_3221gat, id_3157gat);
nor ( id_3280gat, id_3224gat, id_3162gat);
nor ( id_3284gat, id_3227gat, id_3167gat);
nor ( id_3288gat, id_3230gat, id_3172gat);
nor ( id_3292gat, id_3233gat, id_3177gat);
nor ( id_3296gat, id_3236gat, id_3182gat);
nor ( id_3300gat, id_3190gat, id_3239gat);
nor ( id_3301gat, id_3239gat, id_3187gat);
nor ( id_3302gat, id_3243gat, id_3244gat);
nor ( id_3305gat, id_3245gat, id_1092gat);
nor ( id_3309gat, id_3199gat, id_3248gat);
nor ( id_3310gat, id_3248gat, id_1140gat);
nor ( id_3311gat, id_3070gat, id_3248gat);
nor ( id_3314gat, id_3252gat, id_3253gat);
nor ( id_3317gat, id_3257gat, id_3254gat);
nor ( id_3321gat, id_1284gat, id_3260gat);
nor ( id_3322gat, id_3260gat, id_3208gat);
nor ( id_3323gat, id_3212gat, id_3264gat);
nor ( id_3324gat, id_3264gat, id_3142gat);
nor ( id_3325gat, id_3215gat, id_3268gat);
nor ( id_3326gat, id_3268gat, id_3147gat);
nor ( id_3327gat, id_3218gat, id_3272gat);
nor ( id_3328gat, id_3272gat, id_3152gat);
nor ( id_3329gat, id_3221gat, id_3276gat);
nor ( id_3330gat, id_3276gat, id_3157gat);
nor ( id_3331gat, id_3224gat, id_3280gat);
nor ( id_3332gat, id_3280gat, id_3162gat);
nor ( id_3333gat, id_3227gat, id_3284gat);
nor ( id_3334gat, id_3284gat, id_3167gat);
nor ( id_3335gat, id_3230gat, id_3288gat);
nor ( id_3336gat, id_3288gat, id_3172gat);
nor ( id_3337gat, id_3233gat, id_3292gat);
nor ( id_3338gat, id_3292gat, id_3177gat);
nor ( id_3339gat, id_3236gat, id_3296gat);
nor ( id_3340gat, id_3296gat, id_3182gat);
nor ( id_3341gat, id_3300gat, id_3301gat);
nor ( id_3344gat, id_3302gat, id_1044gat);
nor ( id_3348gat, id_3245gat, id_3305gat);
nor ( id_3349gat, id_3305gat, id_1092gat);
nor ( id_3350gat, id_3127gat, id_3305gat);
nor ( id_3353gat, id_3309gat, id_3310gat);
nor ( id_3356gat, id_3314gat, id_3311gat);
nor ( id_3360gat, id_3257gat, id_3317gat);
nor ( id_3361gat, id_3317gat, id_3254gat);
nor ( id_3362gat, id_3321gat, id_3322gat);
nor ( id_3365gat, id_3323gat, id_3324gat);
nor ( id_3368gat, id_3325gat, id_3326gat);
nor ( id_3371gat, id_3327gat, id_3328gat);
nor ( id_3374gat, id_3329gat, id_3330gat);
nor ( id_3377gat, id_3331gat, id_3332gat);
nor ( id_3380gat, id_3333gat, id_3334gat);
nor ( id_3383gat, id_3335gat, id_3336gat);
nor ( id_3386gat, id_3337gat, id_3338gat);
nor ( id_3389gat, id_3339gat, id_3340gat);
nor ( id_3392gat, id_3341gat, id_996gat);
nor ( id_3396gat, id_3302gat, id_3344gat);
nor ( id_3397gat, id_3344gat, id_1044gat);
nor ( id_3398gat, id_3193gat, id_3344gat);
nor ( id_3401gat, id_3348gat, id_3349gat);
nor ( id_3404gat, id_3353gat, id_3350gat);
nor ( id_3408gat, id_3314gat, id_3356gat);
nor ( id_3409gat, id_3356gat, id_3311gat);
nor ( id_3410gat, id_3360gat, id_3361gat);
nor ( id_3413gat, id_3362gat, id_1239gat);
nor ( id_3417gat, id_3365gat, id_564gat);
nor ( id_3421gat, id_3368gat, id_612gat);
nor ( id_3425gat, id_3371gat, id_660gat);
nor ( id_3429gat, id_3374gat, id_708gat);
nor ( id_3433gat, id_3377gat, id_756gat);
nor ( id_3437gat, id_3380gat, id_804gat);
nor ( id_3441gat, id_3383gat, id_852gat);
nor ( id_3445gat, id_3386gat, id_900gat);
nor ( id_3449gat, id_3389gat, id_948gat);
nor ( id_3453gat, id_3341gat, id_3392gat);
nor ( id_3454gat, id_3392gat, id_996gat);
nor ( id_3455gat, id_3239gat, id_3392gat);
nor ( id_3458gat, id_3396gat, id_3397gat);
nor ( id_3461gat, id_3401gat, id_3398gat);
nor ( id_3465gat, id_3353gat, id_3404gat);
nor ( id_3466gat, id_3404gat, id_3350gat);
nor ( id_3467gat, id_3408gat, id_3409gat);
nor ( id_3470gat, id_3410gat, id_1191gat);
nor ( id_3474gat, id_3362gat, id_3413gat);
nor ( id_3475gat, id_3413gat, id_1239gat);
nor ( id_3476gat, id_3260gat, id_3413gat);
nor ( id_3479gat, id_3365gat, id_3417gat);
nor ( id_3480gat, id_3417gat, id_564gat);
nor ( id_3481gat, id_3264gat, id_3417gat);
nor ( id_3484gat, id_3368gat, id_3421gat);
nor ( id_3485gat, id_3421gat, id_612gat);
nor ( id_3486gat, id_3268gat, id_3421gat);
nor ( id_3489gat, id_3371gat, id_3425gat);
nor ( id_3490gat, id_3425gat, id_660gat);
nor ( id_3491gat, id_3272gat, id_3425gat);
nor ( id_3494gat, id_3374gat, id_3429gat);
nor ( id_3495gat, id_3429gat, id_708gat);
nor ( id_3496gat, id_3276gat, id_3429gat);
nor ( id_3499gat, id_3377gat, id_3433gat);
nor ( id_3500gat, id_3433gat, id_756gat);
nor ( id_3501gat, id_3280gat, id_3433gat);
nor ( id_3504gat, id_3380gat, id_3437gat);
nor ( id_3505gat, id_3437gat, id_804gat);
nor ( id_3506gat, id_3284gat, id_3437gat);
nor ( id_3509gat, id_3383gat, id_3441gat);
nor ( id_3510gat, id_3441gat, id_852gat);
nor ( id_3511gat, id_3288gat, id_3441gat);
nor ( id_3514gat, id_3386gat, id_3445gat);
nor ( id_3515gat, id_3445gat, id_900gat);
nor ( id_3516gat, id_3292gat, id_3445gat);
nor ( id_3519gat, id_3389gat, id_3449gat);
nor ( id_3520gat, id_3449gat, id_948gat);
nor ( id_3521gat, id_3296gat, id_3449gat);
nor ( id_3524gat, id_3453gat, id_3454gat);
nor ( id_3527gat, id_3458gat, id_3455gat);
nor ( id_3531gat, id_3401gat, id_3461gat);
nor ( id_3532gat, id_3461gat, id_3398gat);
nor ( id_3533gat, id_3465gat, id_3466gat);
nor ( id_3536gat, id_3467gat, id_1143gat);
nor ( id_3540gat, id_3410gat, id_3470gat);
nor ( id_3541gat, id_3470gat, id_1191gat);
nor ( id_3542gat, id_3317gat, id_3470gat);
nor ( id_3545gat, id_3474gat, id_3475gat);
nor ( id_3548gat, id_1287gat, id_3476gat);
nor ( id_3552gat, id_3479gat, id_3480gat);
nor ( id_3553gat, id_3484gat, id_3485gat);
nor ( id_3556gat, id_3489gat, id_3490gat);
nor ( id_3559gat, id_3494gat, id_3495gat);
nor ( id_3562gat, id_3499gat, id_3500gat);
nor ( id_3565gat, id_3504gat, id_3505gat);
nor ( id_3568gat, id_3509gat, id_3510gat);
nor ( id_3571gat, id_3514gat, id_3515gat);
nor ( id_3574gat, id_3519gat, id_3520gat);
nor ( id_3577gat, id_3524gat, id_3521gat);
nor ( id_3581gat, id_3458gat, id_3527gat);
nor ( id_3582gat, id_3527gat, id_3455gat);
nor ( id_3583gat, id_3531gat, id_3532gat);
nor ( id_3586gat, id_3533gat, id_1095gat);
nor ( id_3590gat, id_3467gat, id_3536gat);
nor ( id_3591gat, id_3536gat, id_1143gat);
nor ( id_3592gat, id_3356gat, id_3536gat);
nor ( id_3595gat, id_3540gat, id_3541gat);
nor ( id_3598gat, id_3545gat, id_3542gat);
nor ( id_3602gat, id_1287gat, id_3548gat);
nor ( id_3603gat, id_3548gat, id_3476gat);
nor ( id_3604gat, id_3553gat, id_3481gat);
nor ( id_3608gat, id_3556gat, id_3486gat);
nor ( id_3612gat, id_3559gat, id_3491gat);
nor ( id_3616gat, id_3562gat, id_3496gat);
nor ( id_3620gat, id_3565gat, id_3501gat);
nor ( id_3624gat, id_3568gat, id_3506gat);
nor ( id_3628gat, id_3571gat, id_3511gat);
nor ( id_3632gat, id_3574gat, id_3516gat);
nor ( id_3636gat, id_3524gat, id_3577gat);
nor ( id_3637gat, id_3577gat, id_3521gat);
nor ( id_3638gat, id_3581gat, id_3582gat);
nor ( id_3641gat, id_3583gat, id_1047gat);
nor ( id_3645gat, id_3533gat, id_3586gat);
nor ( id_3646gat, id_3586gat, id_1095gat);
nor ( id_3647gat, id_3404gat, id_3586gat);
nor ( id_3650gat, id_3590gat, id_3591gat);
nor ( id_3653gat, id_3595gat, id_3592gat);
nor ( id_3657gat, id_3545gat, id_3598gat);
nor ( id_3658gat, id_3598gat, id_3542gat);
nor ( id_3659gat, id_3602gat, id_3603gat);
nor ( id_3662gat, id_3553gat, id_3604gat);
nor ( id_3663gat, id_3604gat, id_3481gat);
nor ( id_3664gat, id_3556gat, id_3608gat);
nor ( id_3665gat, id_3608gat, id_3486gat);
nor ( id_3666gat, id_3559gat, id_3612gat);
nor ( id_3667gat, id_3612gat, id_3491gat);
nor ( id_3668gat, id_3562gat, id_3616gat);
nor ( id_3669gat, id_3616gat, id_3496gat);
nor ( id_3670gat, id_3565gat, id_3620gat);
nor ( id_3671gat, id_3620gat, id_3501gat);
nor ( id_3672gat, id_3568gat, id_3624gat);
nor ( id_3673gat, id_3624gat, id_3506gat);
nor ( id_3674gat, id_3571gat, id_3628gat);
nor ( id_3675gat, id_3628gat, id_3511gat);
nor ( id_3676gat, id_3574gat, id_3632gat);
nor ( id_3677gat, id_3632gat, id_3516gat);
nor ( id_3678gat, id_3636gat, id_3637gat);
nor ( id_3681gat, id_3638gat, id_999gat);
nor ( id_3685gat, id_3583gat, id_3641gat);
nor ( id_3686gat, id_3641gat, id_1047gat);
nor ( id_3687gat, id_3461gat, id_3641gat);
nor ( id_3690gat, id_3645gat, id_3646gat);
nor ( id_3693gat, id_3650gat, id_3647gat);
nor ( id_3697gat, id_3595gat, id_3653gat);
nor ( id_3698gat, id_3653gat, id_3592gat);
nor ( id_3699gat, id_3657gat, id_3658gat);
nor ( id_3702gat, id_3659gat, id_1242gat);
nor ( id_3706gat, id_3662gat, id_3663gat);
nor ( id_3709gat, id_3664gat, id_3665gat);
nor ( id_3712gat, id_3666gat, id_3667gat);
nor ( id_3715gat, id_3668gat, id_3669gat);
nor ( id_3718gat, id_3670gat, id_3671gat);
nor ( id_3721gat, id_3672gat, id_3673gat);
nor ( id_3724gat, id_3674gat, id_3675gat);
nor ( id_3727gat, id_3676gat, id_3677gat);
nor ( id_3730gat, id_3678gat, id_951gat);
nor ( id_3734gat, id_3638gat, id_3681gat);
nor ( id_3735gat, id_3681gat, id_999gat);
nor ( id_3736gat, id_3527gat, id_3681gat);
nor ( id_3739gat, id_3685gat, id_3686gat);
nor ( id_3742gat, id_3690gat, id_3687gat);
nor ( id_3746gat, id_3650gat, id_3693gat);
nor ( id_3747gat, id_3693gat, id_3647gat);
nor ( id_3748gat, id_3697gat, id_3698gat);
nor ( id_3751gat, id_3699gat, id_1194gat);
nor ( id_3755gat, id_3659gat, id_3702gat);
nor ( id_3756gat, id_3702gat, id_1242gat);
nor ( id_3757gat, id_3548gat, id_3702gat);
nor ( id_3760gat, id_3706gat, id_567gat);
nor ( id_3764gat, id_3709gat, id_615gat);
nor ( id_3768gat, id_3712gat, id_663gat);
nor ( id_3772gat, id_3715gat, id_711gat);
nor ( id_3776gat, id_3718gat, id_759gat);
nor ( id_3780gat, id_3721gat, id_807gat);
nor ( id_3784gat, id_3724gat, id_855gat);
nor ( id_3788gat, id_3727gat, id_903gat);
nor ( id_3792gat, id_3678gat, id_3730gat);
nor ( id_3793gat, id_3730gat, id_951gat);
nor ( id_3794gat, id_3577gat, id_3730gat);
nor ( id_3797gat, id_3734gat, id_3735gat);
nor ( id_3800gat, id_3739gat, id_3736gat);
nor ( id_3804gat, id_3690gat, id_3742gat);
nor ( id_3805gat, id_3742gat, id_3687gat);
nor ( id_3806gat, id_3746gat, id_3747gat);
nor ( id_3809gat, id_3748gat, id_1146gat);
nor ( id_3813gat, id_3699gat, id_3751gat);
nor ( id_3814gat, id_3751gat, id_1194gat);
nor ( id_3815gat, id_3598gat, id_3751gat);
nor ( id_3818gat, id_3755gat, id_3756gat);
nor ( id_3821gat, id_1290gat, id_3757gat);
nor ( id_3825gat, id_3706gat, id_3760gat);
nor ( id_3826gat, id_3760gat, id_567gat);
nor ( id_3827gat, id_3604gat, id_3760gat);
nor ( id_3830gat, id_3709gat, id_3764gat);
nor ( id_3831gat, id_3764gat, id_615gat);
nor ( id_3832gat, id_3608gat, id_3764gat);
nor ( id_3835gat, id_3712gat, id_3768gat);
nor ( id_3836gat, id_3768gat, id_663gat);
nor ( id_3837gat, id_3612gat, id_3768gat);
nor ( id_3840gat, id_3715gat, id_3772gat);
nor ( id_3841gat, id_3772gat, id_711gat);
nor ( id_3842gat, id_3616gat, id_3772gat);
nor ( id_3845gat, id_3718gat, id_3776gat);
nor ( id_3846gat, id_3776gat, id_759gat);
nor ( id_3847gat, id_3620gat, id_3776gat);
nor ( id_3850gat, id_3721gat, id_3780gat);
nor ( id_3851gat, id_3780gat, id_807gat);
nor ( id_3852gat, id_3624gat, id_3780gat);
nor ( id_3855gat, id_3724gat, id_3784gat);
nor ( id_3856gat, id_3784gat, id_855gat);
nor ( id_3857gat, id_3628gat, id_3784gat);
nor ( id_3860gat, id_3727gat, id_3788gat);
nor ( id_3861gat, id_3788gat, id_903gat);
nor ( id_3862gat, id_3632gat, id_3788gat);
nor ( id_3865gat, id_3792gat, id_3793gat);
nor ( id_3868gat, id_3797gat, id_3794gat);
nor ( id_3872gat, id_3739gat, id_3800gat);
nor ( id_3873gat, id_3800gat, id_3736gat);
nor ( id_3874gat, id_3804gat, id_3805gat);
nor ( id_3877gat, id_3806gat, id_1098gat);
nor ( id_3881gat, id_3748gat, id_3809gat);
nor ( id_3882gat, id_3809gat, id_1146gat);
nor ( id_3883gat, id_3653gat, id_3809gat);
nor ( id_3886gat, id_3813gat, id_3814gat);
nor ( id_3889gat, id_3818gat, id_3815gat);
nor ( id_3893gat, id_1290gat, id_3821gat);
nor ( id_3894gat, id_3821gat, id_3757gat);
nor ( id_3895gat, id_3825gat, id_3826gat);
nor ( id_3896gat, id_3830gat, id_3831gat);
nor ( id_3899gat, id_3835gat, id_3836gat);
nor ( id_3902gat, id_3840gat, id_3841gat);
nor ( id_3905gat, id_3845gat, id_3846gat);
nor ( id_3908gat, id_3850gat, id_3851gat);
nor ( id_3911gat, id_3855gat, id_3856gat);
nor ( id_3914gat, id_3860gat, id_3861gat);
nor ( id_3917gat, id_3865gat, id_3862gat);
nor ( id_3921gat, id_3797gat, id_3868gat);
nor ( id_3922gat, id_3868gat, id_3794gat);
nor ( id_3923gat, id_3872gat, id_3873gat);
nor ( id_3926gat, id_3874gat, id_1050gat);
nor ( id_3930gat, id_3806gat, id_3877gat);
nor ( id_3931gat, id_3877gat, id_1098gat);
nor ( id_3932gat, id_3693gat, id_3877gat);
nor ( id_3935gat, id_3881gat, id_3882gat);
nor ( id_3938gat, id_3886gat, id_3883gat);
nor ( id_3942gat, id_3818gat, id_3889gat);
nor ( id_3943gat, id_3889gat, id_3815gat);
nor ( id_3944gat, id_3893gat, id_3894gat);
nor ( id_3947gat, id_3896gat, id_3827gat);
nor ( id_3951gat, id_3899gat, id_3832gat);
nor ( id_3955gat, id_3902gat, id_3837gat);
nor ( id_3959gat, id_3905gat, id_3842gat);
nor ( id_3963gat, id_3908gat, id_3847gat);
nor ( id_3967gat, id_3911gat, id_3852gat);
nor ( id_3971gat, id_3914gat, id_3857gat);
nor ( id_3975gat, id_3865gat, id_3917gat);
nor ( id_3976gat, id_3917gat, id_3862gat);
nor ( id_3977gat, id_3921gat, id_3922gat);
nor ( id_3980gat, id_3923gat, id_1002gat);
nor ( id_3984gat, id_3874gat, id_3926gat);
nor ( id_3985gat, id_3926gat, id_1050gat);
nor ( id_3986gat, id_3742gat, id_3926gat);
nor ( id_3989gat, id_3930gat, id_3931gat);
nor ( id_3992gat, id_3935gat, id_3932gat);
nor ( id_3996gat, id_3886gat, id_3938gat);
nor ( id_3997gat, id_3938gat, id_3883gat);
nor ( id_3998gat, id_3942gat, id_3943gat);
nor ( id_4001gat, id_3944gat, id_1245gat);
nor ( id_4005gat, id_3896gat, id_3947gat);
nor ( id_4006gat, id_3947gat, id_3827gat);
nor ( id_4007gat, id_3899gat, id_3951gat);
nor ( id_4008gat, id_3951gat, id_3832gat);
nor ( id_4009gat, id_3902gat, id_3955gat);
nor ( id_4010gat, id_3955gat, id_3837gat);
nor ( id_4011gat, id_3905gat, id_3959gat);
nor ( id_4012gat, id_3959gat, id_3842gat);
nor ( id_4013gat, id_3908gat, id_3963gat);
nor ( id_4014gat, id_3963gat, id_3847gat);
nor ( id_4015gat, id_3911gat, id_3967gat);
nor ( id_4016gat, id_3967gat, id_3852gat);
nor ( id_4017gat, id_3914gat, id_3971gat);
nor ( id_4018gat, id_3971gat, id_3857gat);
nor ( id_4019gat, id_3975gat, id_3976gat);
nor ( id_4022gat, id_3977gat, id_954gat);
nor ( id_4026gat, id_3923gat, id_3980gat);
nor ( id_4027gat, id_3980gat, id_1002gat);
nor ( id_4028gat, id_3800gat, id_3980gat);
nor ( id_4031gat, id_3984gat, id_3985gat);
nor ( id_4034gat, id_3989gat, id_3986gat);
nor ( id_4038gat, id_3935gat, id_3992gat);
nor ( id_4039gat, id_3992gat, id_3932gat);
nor ( id_4040gat, id_3996gat, id_3997gat);
nor ( id_4043gat, id_3998gat, id_1197gat);
nor ( id_4047gat, id_3944gat, id_4001gat);
nor ( id_4048gat, id_4001gat, id_1245gat);
nor ( id_4049gat, id_3821gat, id_4001gat);
nor ( id_4052gat, id_4005gat, id_4006gat);
nor ( id_4055gat, id_4007gat, id_4008gat);
nor ( id_4058gat, id_4009gat, id_4010gat);
nor ( id_4061gat, id_4011gat, id_4012gat);
nor ( id_4064gat, id_4013gat, id_4014gat);
nor ( id_4067gat, id_4015gat, id_4016gat);
nor ( id_4070gat, id_4017gat, id_4018gat);
nor ( id_4073gat, id_4019gat, id_906gat);
nor ( id_4077gat, id_3977gat, id_4022gat);
nor ( id_4078gat, id_4022gat, id_954gat);
nor ( id_4079gat, id_3868gat, id_4022gat);
nor ( id_4082gat, id_4026gat, id_4027gat);
nor ( id_4085gat, id_4031gat, id_4028gat);
nor ( id_4089gat, id_3989gat, id_4034gat);
nor ( id_4090gat, id_4034gat, id_3986gat);
nor ( id_4091gat, id_4038gat, id_4039gat);
nor ( id_4094gat, id_4040gat, id_1149gat);
nor ( id_4098gat, id_3998gat, id_4043gat);
nor ( id_4099gat, id_4043gat, id_1197gat);
nor ( id_4100gat, id_3889gat, id_4043gat);
nor ( id_4103gat, id_4047gat, id_4048gat);
nor ( id_4106gat, id_1293gat, id_4049gat);
nor ( id_4110gat, id_4052gat, id_570gat);
nor ( id_4114gat, id_4055gat, id_618gat);
nor ( id_4118gat, id_4058gat, id_666gat);
nor ( id_4122gat, id_4061gat, id_714gat);
nor ( id_4126gat, id_4064gat, id_762gat);
nor ( id_4130gat, id_4067gat, id_810gat);
nor ( id_4134gat, id_4070gat, id_858gat);
nor ( id_4138gat, id_4019gat, id_4073gat);
nor ( id_4139gat, id_4073gat, id_906gat);
nor ( id_4140gat, id_3917gat, id_4073gat);
nor ( id_4143gat, id_4077gat, id_4078gat);
nor ( id_4146gat, id_4082gat, id_4079gat);
nor ( id_4150gat, id_4031gat, id_4085gat);
nor ( id_4151gat, id_4085gat, id_4028gat);
nor ( id_4152gat, id_4089gat, id_4090gat);
nor ( id_4155gat, id_4091gat, id_1101gat);
nor ( id_4159gat, id_4040gat, id_4094gat);
nor ( id_4160gat, id_4094gat, id_1149gat);
nor ( id_4161gat, id_3938gat, id_4094gat);
nor ( id_4164gat, id_4098gat, id_4099gat);
nor ( id_4167gat, id_4103gat, id_4100gat);
nor ( id_4171gat, id_1293gat, id_4106gat);
nor ( id_4172gat, id_4106gat, id_4049gat);
nor ( id_4173gat, id_4052gat, id_4110gat);
nor ( id_4174gat, id_4110gat, id_570gat);
nor ( id_4175gat, id_3947gat, id_4110gat);
nor ( id_4178gat, id_4055gat, id_4114gat);
nor ( id_4179gat, id_4114gat, id_618gat);
nor ( id_4180gat, id_3951gat, id_4114gat);
nor ( id_4183gat, id_4058gat, id_4118gat);
nor ( id_4184gat, id_4118gat, id_666gat);
nor ( id_4185gat, id_3955gat, id_4118gat);
nor ( id_4188gat, id_4061gat, id_4122gat);
nor ( id_4189gat, id_4122gat, id_714gat);
nor ( id_4190gat, id_3959gat, id_4122gat);
nor ( id_4193gat, id_4064gat, id_4126gat);
nor ( id_4194gat, id_4126gat, id_762gat);
nor ( id_4195gat, id_3963gat, id_4126gat);
nor ( id_4198gat, id_4067gat, id_4130gat);
nor ( id_4199gat, id_4130gat, id_810gat);
nor ( id_4200gat, id_3967gat, id_4130gat);
nor ( id_4203gat, id_4070gat, id_4134gat);
nor ( id_4204gat, id_4134gat, id_858gat);
nor ( id_4205gat, id_3971gat, id_4134gat);
nor ( id_4208gat, id_4138gat, id_4139gat);
nor ( id_4211gat, id_4143gat, id_4140gat);
nor ( id_4215gat, id_4082gat, id_4146gat);
nor ( id_4216gat, id_4146gat, id_4079gat);
nor ( id_4217gat, id_4150gat, id_4151gat);
nor ( id_4220gat, id_4152gat, id_1053gat);
nor ( id_4224gat, id_4091gat, id_4155gat);
nor ( id_4225gat, id_4155gat, id_1101gat);
nor ( id_4226gat, id_3992gat, id_4155gat);
nor ( id_4229gat, id_4159gat, id_4160gat);
nor ( id_4232gat, id_4164gat, id_4161gat);
nor ( id_4236gat, id_4103gat, id_4167gat);
nor ( id_4237gat, id_4167gat, id_4100gat);
nor ( id_4238gat, id_4171gat, id_4172gat);
nor ( id_4241gat, id_4173gat, id_4174gat);
nor ( id_4242gat, id_4178gat, id_4179gat);
nor ( id_4245gat, id_4183gat, id_4184gat);
nor ( id_4248gat, id_4188gat, id_4189gat);
nor ( id_4251gat, id_4193gat, id_4194gat);
nor ( id_4254gat, id_4198gat, id_4199gat);
nor ( id_4257gat, id_4203gat, id_4204gat);
nor ( id_4260gat, id_4208gat, id_4205gat);
nor ( id_4264gat, id_4143gat, id_4211gat);
nor ( id_4265gat, id_4211gat, id_4140gat);
nor ( id_4266gat, id_4215gat, id_4216gat);
nor ( id_4269gat, id_4217gat, id_1005gat);
nor ( id_4273gat, id_4152gat, id_4220gat);
nor ( id_4274gat, id_4220gat, id_1053gat);
nor ( id_4275gat, id_4034gat, id_4220gat);
nor ( id_4278gat, id_4224gat, id_4225gat);
nor ( id_4281gat, id_4229gat, id_4226gat);
nor ( id_4285gat, id_4164gat, id_4232gat);
nor ( id_4286gat, id_4232gat, id_4161gat);
nor ( id_4287gat, id_4236gat, id_4237gat);
nor ( id_4290gat, id_4238gat, id_1248gat);
nor ( id_4294gat, id_4242gat, id_4175gat);
nor ( id_4298gat, id_4245gat, id_4180gat);
nor ( id_4302gat, id_4248gat, id_4185gat);
nor ( id_4306gat, id_4251gat, id_4190gat);
nor ( id_4310gat, id_4254gat, id_4195gat);
nor ( id_4314gat, id_4257gat, id_4200gat);
nor ( id_4318gat, id_4208gat, id_4260gat);
nor ( id_4319gat, id_4260gat, id_4205gat);
nor ( id_4320gat, id_4264gat, id_4265gat);
nor ( id_4323gat, id_4266gat, id_957gat);
nor ( id_4327gat, id_4217gat, id_4269gat);
nor ( id_4328gat, id_4269gat, id_1005gat);
nor ( id_4329gat, id_4085gat, id_4269gat);
nor ( id_4332gat, id_4273gat, id_4274gat);
nor ( id_4335gat, id_4278gat, id_4275gat);
nor ( id_4339gat, id_4229gat, id_4281gat);
nor ( id_4340gat, id_4281gat, id_4226gat);
nor ( id_4341gat, id_4285gat, id_4286gat);
nor ( id_4344gat, id_4287gat, id_1200gat);
nor ( id_4348gat, id_4238gat, id_4290gat);
nor ( id_4349gat, id_4290gat, id_1248gat);
nor ( id_4350gat, id_4106gat, id_4290gat);
nor ( id_4353gat, id_4242gat, id_4294gat);
nor ( id_4354gat, id_4294gat, id_4175gat);
nor ( id_4355gat, id_4245gat, id_4298gat);
nor ( id_4356gat, id_4298gat, id_4180gat);
nor ( id_4357gat, id_4248gat, id_4302gat);
nor ( id_4358gat, id_4302gat, id_4185gat);
nor ( id_4359gat, id_4251gat, id_4306gat);
nor ( id_4360gat, id_4306gat, id_4190gat);
nor ( id_4361gat, id_4254gat, id_4310gat);
nor ( id_4362gat, id_4310gat, id_4195gat);
nor ( id_4363gat, id_4257gat, id_4314gat);
nor ( id_4364gat, id_4314gat, id_4200gat);
nor ( id_4365gat, id_4318gat, id_4319gat);
nor ( id_4368gat, id_4320gat, id_909gat);
nor ( id_4372gat, id_4266gat, id_4323gat);
nor ( id_4373gat, id_4323gat, id_957gat);
nor ( id_4374gat, id_4146gat, id_4323gat);
nor ( id_4377gat, id_4327gat, id_4328gat);
nor ( id_4380gat, id_4332gat, id_4329gat);
nor ( id_4384gat, id_4278gat, id_4335gat);
nor ( id_4385gat, id_4335gat, id_4275gat);
nor ( id_4386gat, id_4339gat, id_4340gat);
nor ( id_4389gat, id_4341gat, id_1152gat);
nor ( id_4393gat, id_4287gat, id_4344gat);
nor ( id_4394gat, id_4344gat, id_1200gat);
nor ( id_4395gat, id_4167gat, id_4344gat);
nor ( id_4398gat, id_4348gat, id_4349gat);
nor ( id_4401gat, id_1296gat, id_4350gat);
nor ( id_4405gat, id_4353gat, id_4354gat);
nor ( id_4408gat, id_4355gat, id_4356gat);
nor ( id_4411gat, id_4357gat, id_4358gat);
nor ( id_4414gat, id_4359gat, id_4360gat);
nor ( id_4417gat, id_4361gat, id_4362gat);
nor ( id_4420gat, id_4363gat, id_4364gat);
nor ( id_4423gat, id_4365gat, id_861gat);
nor ( id_4427gat, id_4320gat, id_4368gat);
nor ( id_4428gat, id_4368gat, id_909gat);
nor ( id_4429gat, id_4211gat, id_4368gat);
nor ( id_4432gat, id_4372gat, id_4373gat);
nor ( id_4435gat, id_4377gat, id_4374gat);
nor ( id_4439gat, id_4332gat, id_4380gat);
nor ( id_4440gat, id_4380gat, id_4329gat);
nor ( id_4441gat, id_4384gat, id_4385gat);
nor ( id_4444gat, id_4386gat, id_1104gat);
nor ( id_4448gat, id_4341gat, id_4389gat);
nor ( id_4449gat, id_4389gat, id_1152gat);
nor ( id_4450gat, id_4232gat, id_4389gat);
nor ( id_4453gat, id_4393gat, id_4394gat);
nor ( id_4456gat, id_4398gat, id_4395gat);
nor ( id_4460gat, id_1296gat, id_4401gat);
nor ( id_4461gat, id_4401gat, id_4350gat);
nor ( id_4462gat, id_4405gat, id_573gat);
nor ( id_4466gat, id_4408gat, id_621gat);
nor ( id_4470gat, id_4411gat, id_669gat);
nor ( id_4474gat, id_4414gat, id_717gat);
nor ( id_4478gat, id_4417gat, id_765gat);
nor ( id_4482gat, id_4420gat, id_813gat);
nor ( id_4486gat, id_4365gat, id_4423gat);
nor ( id_4487gat, id_4423gat, id_861gat);
nor ( id_4488gat, id_4260gat, id_4423gat);
nor ( id_4491gat, id_4427gat, id_4428gat);
nor ( id_4494gat, id_4432gat, id_4429gat);
nor ( id_4498gat, id_4377gat, id_4435gat);
nor ( id_4499gat, id_4435gat, id_4374gat);
nor ( id_4500gat, id_4439gat, id_4440gat);
nor ( id_4503gat, id_4441gat, id_1056gat);
nor ( id_4507gat, id_4386gat, id_4444gat);
nor ( id_4508gat, id_4444gat, id_1104gat);
nor ( id_4509gat, id_4281gat, id_4444gat);
nor ( id_4512gat, id_4448gat, id_4449gat);
nor ( id_4515gat, id_4453gat, id_4450gat);
nor ( id_4519gat, id_4398gat, id_4456gat);
nor ( id_4520gat, id_4456gat, id_4395gat);
nor ( id_4521gat, id_4460gat, id_4461gat);
nor ( id_4524gat, id_4405gat, id_4462gat);
nor ( id_4525gat, id_4462gat, id_573gat);
nor ( id_4526gat, id_4294gat, id_4462gat);
nor ( id_4529gat, id_4408gat, id_4466gat);
nor ( id_4530gat, id_4466gat, id_621gat);
nor ( id_4531gat, id_4298gat, id_4466gat);
nor ( id_4534gat, id_4411gat, id_4470gat);
nor ( id_4535gat, id_4470gat, id_669gat);
nor ( id_4536gat, id_4302gat, id_4470gat);
nor ( id_4539gat, id_4414gat, id_4474gat);
nor ( id_4540gat, id_4474gat, id_717gat);
nor ( id_4541gat, id_4306gat, id_4474gat);
nor ( id_4544gat, id_4417gat, id_4478gat);
nor ( id_4545gat, id_4478gat, id_765gat);
nor ( id_4546gat, id_4310gat, id_4478gat);
nor ( id_4549gat, id_4420gat, id_4482gat);
nor ( id_4550gat, id_4482gat, id_813gat);
nor ( id_4551gat, id_4314gat, id_4482gat);
nor ( id_4554gat, id_4486gat, id_4487gat);
nor ( id_4557gat, id_4491gat, id_4488gat);
nor ( id_4561gat, id_4432gat, id_4494gat);
nor ( id_4562gat, id_4494gat, id_4429gat);
nor ( id_4563gat, id_4498gat, id_4499gat);
nor ( id_4566gat, id_4500gat, id_1008gat);
nor ( id_4570gat, id_4441gat, id_4503gat);
nor ( id_4571gat, id_4503gat, id_1056gat);
nor ( id_4572gat, id_4335gat, id_4503gat);
nor ( id_4575gat, id_4507gat, id_4508gat);
nor ( id_4578gat, id_4512gat, id_4509gat);
nor ( id_4582gat, id_4453gat, id_4515gat);
nor ( id_4583gat, id_4515gat, id_4450gat);
nor ( id_4584gat, id_4519gat, id_4520gat);
nor ( id_4587gat, id_4521gat, id_1251gat);
nor ( id_4591gat, id_4524gat, id_4525gat);
nor ( id_4592gat, id_4529gat, id_4530gat);
nor ( id_4595gat, id_4534gat, id_4535gat);
nor ( id_4598gat, id_4539gat, id_4540gat);
nor ( id_4601gat, id_4544gat, id_4545gat);
nor ( id_4604gat, id_4549gat, id_4550gat);
nor ( id_4607gat, id_4554gat, id_4551gat);
nor ( id_4611gat, id_4491gat, id_4557gat);
nor ( id_4612gat, id_4557gat, id_4488gat);
nor ( id_4613gat, id_4561gat, id_4562gat);
nor ( id_4616gat, id_4563gat, id_960gat);
nor ( id_4620gat, id_4500gat, id_4566gat);
nor ( id_4621gat, id_4566gat, id_1008gat);
nor ( id_4622gat, id_4380gat, id_4566gat);
nor ( id_4625gat, id_4570gat, id_4571gat);
nor ( id_4628gat, id_4575gat, id_4572gat);
nor ( id_4632gat, id_4512gat, id_4578gat);
nor ( id_4633gat, id_4578gat, id_4509gat);
nor ( id_4634gat, id_4582gat, id_4583gat);
nor ( id_4637gat, id_4584gat, id_1203gat);
nor ( id_4641gat, id_4521gat, id_4587gat);
nor ( id_4642gat, id_4587gat, id_1251gat);
nor ( id_4643gat, id_4401gat, id_4587gat);
nor ( id_4646gat, id_4592gat, id_4526gat);
nor ( id_4650gat, id_4595gat, id_4531gat);
nor ( id_4654gat, id_4598gat, id_4536gat);
nor ( id_4658gat, id_4601gat, id_4541gat);
nor ( id_4662gat, id_4604gat, id_4546gat);
nor ( id_4666gat, id_4554gat, id_4607gat);
nor ( id_4667gat, id_4607gat, id_4551gat);
nor ( id_4668gat, id_4611gat, id_4612gat);
nor ( id_4671gat, id_4613gat, id_912gat);
nor ( id_4675gat, id_4563gat, id_4616gat);
nor ( id_4676gat, id_4616gat, id_960gat);
nor ( id_4677gat, id_4435gat, id_4616gat);
nor ( id_4680gat, id_4620gat, id_4621gat);
nor ( id_4683gat, id_4625gat, id_4622gat);
nor ( id_4687gat, id_4575gat, id_4628gat);
nor ( id_4688gat, id_4628gat, id_4572gat);
nor ( id_4689gat, id_4632gat, id_4633gat);
nor ( id_4692gat, id_4634gat, id_1155gat);
nor ( id_4696gat, id_4584gat, id_4637gat);
nor ( id_4697gat, id_4637gat, id_1203gat);
nor ( id_4698gat, id_4456gat, id_4637gat);
nor ( id_4701gat, id_4641gat, id_4642gat);
nor ( id_4704gat, id_1299gat, id_4643gat);
nor ( id_4708gat, id_4592gat, id_4646gat);
nor ( id_4709gat, id_4646gat, id_4526gat);
nor ( id_4710gat, id_4595gat, id_4650gat);
nor ( id_4711gat, id_4650gat, id_4531gat);
nor ( id_4712gat, id_4598gat, id_4654gat);
nor ( id_4713gat, id_4654gat, id_4536gat);
nor ( id_4714gat, id_4601gat, id_4658gat);
nor ( id_4715gat, id_4658gat, id_4541gat);
nor ( id_4716gat, id_4604gat, id_4662gat);
nor ( id_4717gat, id_4662gat, id_4546gat);
nor ( id_4718gat, id_4666gat, id_4667gat);
nor ( id_4721gat, id_4668gat, id_864gat);
nor ( id_4725gat, id_4613gat, id_4671gat);
nor ( id_4726gat, id_4671gat, id_912gat);
nor ( id_4727gat, id_4494gat, id_4671gat);
nor ( id_4730gat, id_4675gat, id_4676gat);
nor ( id_4733gat, id_4680gat, id_4677gat);
nor ( id_4737gat, id_4625gat, id_4683gat);
nor ( id_4738gat, id_4683gat, id_4622gat);
nor ( id_4739gat, id_4687gat, id_4688gat);
nor ( id_4742gat, id_4689gat, id_1107gat);
nor ( id_4746gat, id_4634gat, id_4692gat);
nor ( id_4747gat, id_4692gat, id_1155gat);
nor ( id_4748gat, id_4515gat, id_4692gat);
nor ( id_4751gat, id_4696gat, id_4697gat);
nor ( id_4754gat, id_4701gat, id_4698gat);
nor ( id_4758gat, id_1299gat, id_4704gat);
nor ( id_4759gat, id_4704gat, id_4643gat);
nor ( id_4760gat, id_4708gat, id_4709gat);
nor ( id_4763gat, id_4710gat, id_4711gat);
nor ( id_4766gat, id_4712gat, id_4713gat);
nor ( id_4769gat, id_4714gat, id_4715gat);
nor ( id_4772gat, id_4716gat, id_4717gat);
nor ( id_4775gat, id_4718gat, id_816gat);
nor ( id_4779gat, id_4668gat, id_4721gat);
nor ( id_4780gat, id_4721gat, id_864gat);
nor ( id_4781gat, id_4557gat, id_4721gat);
nor ( id_4784gat, id_4725gat, id_4726gat);
nor ( id_4787gat, id_4730gat, id_4727gat);
nor ( id_4791gat, id_4680gat, id_4733gat);
nor ( id_4792gat, id_4733gat, id_4677gat);
nor ( id_4793gat, id_4737gat, id_4738gat);
nor ( id_4796gat, id_4739gat, id_1059gat);
nor ( id_4800gat, id_4689gat, id_4742gat);
nor ( id_4801gat, id_4742gat, id_1107gat);
nor ( id_4802gat, id_4578gat, id_4742gat);
nor ( id_4805gat, id_4746gat, id_4747gat);
nor ( id_4808gat, id_4751gat, id_4748gat);
nor ( id_4812gat, id_4701gat, id_4754gat);
nor ( id_4813gat, id_4754gat, id_4698gat);
nor ( id_4814gat, id_4758gat, id_4759gat);
nor ( id_4817gat, id_4760gat, id_576gat);
nor ( id_4821gat, id_4763gat, id_624gat);
nor ( id_4825gat, id_4766gat, id_672gat);
nor ( id_4829gat, id_4769gat, id_720gat);
nor ( id_4833gat, id_4772gat, id_768gat);
nor ( id_4837gat, id_4718gat, id_4775gat);
nor ( id_4838gat, id_4775gat, id_816gat);
nor ( id_4839gat, id_4607gat, id_4775gat);
nor ( id_4842gat, id_4779gat, id_4780gat);
nor ( id_4845gat, id_4784gat, id_4781gat);
nor ( id_4849gat, id_4730gat, id_4787gat);
nor ( id_4850gat, id_4787gat, id_4727gat);
nor ( id_4851gat, id_4791gat, id_4792gat);
nor ( id_4854gat, id_4793gat, id_1011gat);
nor ( id_4858gat, id_4739gat, id_4796gat);
nor ( id_4859gat, id_4796gat, id_1059gat);
nor ( id_4860gat, id_4628gat, id_4796gat);
nor ( id_4863gat, id_4800gat, id_4801gat);
nor ( id_4866gat, id_4805gat, id_4802gat);
nor ( id_4870gat, id_4751gat, id_4808gat);
nor ( id_4871gat, id_4808gat, id_4748gat);
nor ( id_4872gat, id_4812gat, id_4813gat);
nor ( id_4875gat, id_4814gat, id_1254gat);
nor ( id_4879gat, id_4760gat, id_4817gat);
nor ( id_4880gat, id_4817gat, id_576gat);
nor ( id_4881gat, id_4646gat, id_4817gat);
nor ( id_4884gat, id_4763gat, id_4821gat);
nor ( id_4885gat, id_4821gat, id_624gat);
nor ( id_4886gat, id_4650gat, id_4821gat);
nor ( id_4889gat, id_4766gat, id_4825gat);
nor ( id_4890gat, id_4825gat, id_672gat);
nor ( id_4891gat, id_4654gat, id_4825gat);
nor ( id_4894gat, id_4769gat, id_4829gat);
nor ( id_4895gat, id_4829gat, id_720gat);
nor ( id_4896gat, id_4658gat, id_4829gat);
nor ( id_4899gat, id_4772gat, id_4833gat);
nor ( id_4900gat, id_4833gat, id_768gat);
nor ( id_4901gat, id_4662gat, id_4833gat);
nor ( id_4904gat, id_4837gat, id_4838gat);
nor ( id_4907gat, id_4842gat, id_4839gat);
nor ( id_4911gat, id_4784gat, id_4845gat);
nor ( id_4912gat, id_4845gat, id_4781gat);
nor ( id_4913gat, id_4849gat, id_4850gat);
nor ( id_4916gat, id_4851gat, id_963gat);
nor ( id_4920gat, id_4793gat, id_4854gat);
nor ( id_4921gat, id_4854gat, id_1011gat);
nor ( id_4922gat, id_4683gat, id_4854gat);
nor ( id_4925gat, id_4858gat, id_4859gat);
nor ( id_4928gat, id_4863gat, id_4860gat);
nor ( id_4932gat, id_4805gat, id_4866gat);
nor ( id_4933gat, id_4866gat, id_4802gat);
nor ( id_4934gat, id_4870gat, id_4871gat);
nor ( id_4937gat, id_4872gat, id_1206gat);
nor ( id_4941gat, id_4814gat, id_4875gat);
nor ( id_4942gat, id_4875gat, id_1254gat);
nor ( id_4943gat, id_4704gat, id_4875gat);
nor ( id_4946gat, id_4879gat, id_4880gat);
nor ( id_4947gat, id_4884gat, id_4885gat);
nor ( id_4950gat, id_4889gat, id_4890gat);
nor ( id_4953gat, id_4894gat, id_4895gat);
nor ( id_4956gat, id_4899gat, id_4900gat);
nor ( id_4959gat, id_4904gat, id_4901gat);
nor ( id_4963gat, id_4842gat, id_4907gat);
nor ( id_4964gat, id_4907gat, id_4839gat);
nor ( id_4965gat, id_4911gat, id_4912gat);
nor ( id_4968gat, id_4913gat, id_915gat);
nor ( id_4972gat, id_4851gat, id_4916gat);
nor ( id_4973gat, id_4916gat, id_963gat);
nor ( id_4974gat, id_4733gat, id_4916gat);
nor ( id_4977gat, id_4920gat, id_4921gat);
nor ( id_4980gat, id_4925gat, id_4922gat);
nor ( id_4984gat, id_4863gat, id_4928gat);
nor ( id_4985gat, id_4928gat, id_4860gat);
nor ( id_4986gat, id_4932gat, id_4933gat);
nor ( id_4989gat, id_4934gat, id_1158gat);
nor ( id_4993gat, id_4872gat, id_4937gat);
nor ( id_4994gat, id_4937gat, id_1206gat);
nor ( id_4995gat, id_4754gat, id_4937gat);
nor ( id_4998gat, id_4941gat, id_4942gat);
nor ( id_5001gat, id_1302gat, id_4943gat);
nor ( id_5005gat, id_4947gat, id_4881gat);
nor ( id_5009gat, id_4950gat, id_4886gat);
nor ( id_5013gat, id_4953gat, id_4891gat);
nor ( id_5017gat, id_4956gat, id_4896gat);
nor ( id_5021gat, id_4904gat, id_4959gat);
nor ( id_5022gat, id_4959gat, id_4901gat);
nor ( id_5023gat, id_4963gat, id_4964gat);
nor ( id_5026gat, id_4965gat, id_867gat);
nor ( id_5030gat, id_4913gat, id_4968gat);
nor ( id_5031gat, id_4968gat, id_915gat);
nor ( id_5032gat, id_4787gat, id_4968gat);
nor ( id_5035gat, id_4972gat, id_4973gat);
nor ( id_5038gat, id_4977gat, id_4974gat);
nor ( id_5042gat, id_4925gat, id_4980gat);
nor ( id_5043gat, id_4980gat, id_4922gat);
nor ( id_5044gat, id_4984gat, id_4985gat);
nor ( id_5047gat, id_4986gat, id_1110gat);
nor ( id_5051gat, id_4934gat, id_4989gat);
nor ( id_5052gat, id_4989gat, id_1158gat);
nor ( id_5053gat, id_4808gat, id_4989gat);
nor ( id_5056gat, id_4993gat, id_4994gat);
nor ( id_5059gat, id_4998gat, id_4995gat);
nor ( id_5063gat, id_1302gat, id_5001gat);
nor ( id_5064gat, id_5001gat, id_4943gat);
nor ( id_5065gat, id_4947gat, id_5005gat);
nor ( id_5066gat, id_5005gat, id_4881gat);
nor ( id_5067gat, id_4950gat, id_5009gat);
nor ( id_5068gat, id_5009gat, id_4886gat);
nor ( id_5069gat, id_4953gat, id_5013gat);
nor ( id_5070gat, id_5013gat, id_4891gat);
nor ( id_5071gat, id_4956gat, id_5017gat);
nor ( id_5072gat, id_5017gat, id_4896gat);
nor ( id_5073gat, id_5021gat, id_5022gat);
nor ( id_5076gat, id_5023gat, id_819gat);
nor ( id_5080gat, id_4965gat, id_5026gat);
nor ( id_5081gat, id_5026gat, id_867gat);
nor ( id_5082gat, id_4845gat, id_5026gat);
nor ( id_5085gat, id_5030gat, id_5031gat);
nor ( id_5088gat, id_5035gat, id_5032gat);
nor ( id_5092gat, id_4977gat, id_5038gat);
nor ( id_5093gat, id_5038gat, id_4974gat);
nor ( id_5094gat, id_5042gat, id_5043gat);
nor ( id_5097gat, id_5044gat, id_1062gat);
nor ( id_5101gat, id_4986gat, id_5047gat);
nor ( id_5102gat, id_5047gat, id_1110gat);
nor ( id_5103gat, id_4866gat, id_5047gat);
nor ( id_5106gat, id_5051gat, id_5052gat);
nor ( id_5109gat, id_5056gat, id_5053gat);
nor ( id_5113gat, id_4998gat, id_5059gat);
nor ( id_5114gat, id_5059gat, id_4995gat);
nor ( id_5115gat, id_5063gat, id_5064gat);
nor ( id_5118gat, id_5065gat, id_5066gat);
nor ( id_5121gat, id_5067gat, id_5068gat);
nor ( id_5124gat, id_5069gat, id_5070gat);
nor ( id_5127gat, id_5071gat, id_5072gat);
nor ( id_5130gat, id_5073gat, id_771gat);
nor ( id_5134gat, id_5023gat, id_5076gat);
nor ( id_5135gat, id_5076gat, id_819gat);
nor ( id_5136gat, id_4907gat, id_5076gat);
nor ( id_5139gat, id_5080gat, id_5081gat);
nor ( id_5142gat, id_5085gat, id_5082gat);
nor ( id_5146gat, id_5035gat, id_5088gat);
nor ( id_5147gat, id_5088gat, id_5032gat);
nor ( id_5148gat, id_5092gat, id_5093gat);
nor ( id_5151gat, id_5094gat, id_1014gat);
nor ( id_5155gat, id_5044gat, id_5097gat);
nor ( id_5156gat, id_5097gat, id_1062gat);
nor ( id_5157gat, id_4928gat, id_5097gat);
nor ( id_5160gat, id_5101gat, id_5102gat);
nor ( id_5163gat, id_5106gat, id_5103gat);
nor ( id_5167gat, id_5056gat, id_5109gat);
nor ( id_5168gat, id_5109gat, id_5053gat);
nor ( id_5169gat, id_5113gat, id_5114gat);
nor ( id_5172gat, id_5115gat, id_1257gat);
nor ( id_5176gat, id_5118gat, id_579gat);
nor ( id_5180gat, id_5121gat, id_627gat);
nor ( id_5184gat, id_5124gat, id_675gat);
nor ( id_5188gat, id_5127gat, id_723gat);
nor ( id_5192gat, id_5073gat, id_5130gat);
nor ( id_5193gat, id_5130gat, id_771gat);
nor ( id_5194gat, id_4959gat, id_5130gat);
nor ( id_5197gat, id_5134gat, id_5135gat);
nor ( id_5200gat, id_5139gat, id_5136gat);
nor ( id_5204gat, id_5085gat, id_5142gat);
nor ( id_5205gat, id_5142gat, id_5082gat);
nor ( id_5206gat, id_5146gat, id_5147gat);
nor ( id_5209gat, id_5148gat, id_966gat);
nor ( id_5213gat, id_5094gat, id_5151gat);
nor ( id_5214gat, id_5151gat, id_1014gat);
nor ( id_5215gat, id_4980gat, id_5151gat);
nor ( id_5218gat, id_5155gat, id_5156gat);
nor ( id_5221gat, id_5160gat, id_5157gat);
nor ( id_5225gat, id_5106gat, id_5163gat);
nor ( id_5226gat, id_5163gat, id_5103gat);
nor ( id_5227gat, id_5167gat, id_5168gat);
nor ( id_5230gat, id_5169gat, id_1209gat);
nor ( id_5234gat, id_5115gat, id_5172gat);
nor ( id_5235gat, id_5172gat, id_1257gat);
nor ( id_5236gat, id_5001gat, id_5172gat);
nor ( id_5239gat, id_5118gat, id_5176gat);
nor ( id_5240gat, id_5176gat, id_579gat);
nor ( id_5241gat, id_5005gat, id_5176gat);
nor ( id_5244gat, id_5121gat, id_5180gat);
nor ( id_5245gat, id_5180gat, id_627gat);
nor ( id_5246gat, id_5009gat, id_5180gat);
nor ( id_5249gat, id_5124gat, id_5184gat);
nor ( id_5250gat, id_5184gat, id_675gat);
nor ( id_5251gat, id_5013gat, id_5184gat);
nor ( id_5254gat, id_5127gat, id_5188gat);
nor ( id_5255gat, id_5188gat, id_723gat);
nor ( id_5256gat, id_5017gat, id_5188gat);
nor ( id_5259gat, id_5192gat, id_5193gat);
nor ( id_5262gat, id_5197gat, id_5194gat);
nor ( id_5266gat, id_5139gat, id_5200gat);
nor ( id_5267gat, id_5200gat, id_5136gat);
nor ( id_5268gat, id_5204gat, id_5205gat);
nor ( id_5271gat, id_5206gat, id_918gat);
nor ( id_5275gat, id_5148gat, id_5209gat);
nor ( id_5276gat, id_5209gat, id_966gat);
nor ( id_5277gat, id_5038gat, id_5209gat);
nor ( id_5280gat, id_5213gat, id_5214gat);
nor ( id_5283gat, id_5218gat, id_5215gat);
nor ( id_5287gat, id_5160gat, id_5221gat);
nor ( id_5288gat, id_5221gat, id_5157gat);
nor ( id_5289gat, id_5225gat, id_5226gat);
nor ( id_5292gat, id_5227gat, id_1161gat);
nor ( id_5296gat, id_5169gat, id_5230gat);
nor ( id_5297gat, id_5230gat, id_1209gat);
nor ( id_5298gat, id_5059gat, id_5230gat);
nor ( id_5301gat, id_5234gat, id_5235gat);
nor ( id_5304gat, id_1305gat, id_5236gat);
nor ( id_5308gat, id_5239gat, id_5240gat);
nor ( id_5309gat, id_5244gat, id_5245gat);
nor ( id_5312gat, id_5249gat, id_5250gat);
nor ( id_5315gat, id_5254gat, id_5255gat);
nor ( id_5318gat, id_5259gat, id_5256gat);
nor ( id_5322gat, id_5197gat, id_5262gat);
nor ( id_5323gat, id_5262gat, id_5194gat);
nor ( id_5324gat, id_5266gat, id_5267gat);
nor ( id_5327gat, id_5268gat, id_870gat);
nor ( id_5331gat, id_5206gat, id_5271gat);
nor ( id_5332gat, id_5271gat, id_918gat);
nor ( id_5333gat, id_5088gat, id_5271gat);
nor ( id_5336gat, id_5275gat, id_5276gat);
nor ( id_5339gat, id_5280gat, id_5277gat);
nor ( id_5343gat, id_5218gat, id_5283gat);
nor ( id_5344gat, id_5283gat, id_5215gat);
nor ( id_5345gat, id_5287gat, id_5288gat);
nor ( id_5348gat, id_5289gat, id_1113gat);
nor ( id_5352gat, id_5227gat, id_5292gat);
nor ( id_5353gat, id_5292gat, id_1161gat);
nor ( id_5354gat, id_5109gat, id_5292gat);
nor ( id_5357gat, id_5296gat, id_5297gat);
nor ( id_5360gat, id_5301gat, id_5298gat);
nor ( id_5364gat, id_1305gat, id_5304gat);
nor ( id_5365gat, id_5304gat, id_5236gat);
nor ( id_5366gat, id_5309gat, id_5241gat);
nor ( id_5370gat, id_5312gat, id_5246gat);
nor ( id_5374gat, id_5315gat, id_5251gat);
nor ( id_5378gat, id_5259gat, id_5318gat);
nor ( id_5379gat, id_5318gat, id_5256gat);
nor ( id_5380gat, id_5322gat, id_5323gat);
nor ( id_5383gat, id_5324gat, id_822gat);
nor ( id_5387gat, id_5268gat, id_5327gat);
nor ( id_5388gat, id_5327gat, id_870gat);
nor ( id_5389gat, id_5142gat, id_5327gat);
nor ( id_5392gat, id_5331gat, id_5332gat);
nor ( id_5395gat, id_5336gat, id_5333gat);
nor ( id_5399gat, id_5280gat, id_5339gat);
nor ( id_5400gat, id_5339gat, id_5277gat);
nor ( id_5401gat, id_5343gat, id_5344gat);
nor ( id_5404gat, id_5345gat, id_1065gat);
nor ( id_5408gat, id_5289gat, id_5348gat);
nor ( id_5409gat, id_5348gat, id_1113gat);
nor ( id_5410gat, id_5163gat, id_5348gat);
nor ( id_5413gat, id_5352gat, id_5353gat);
nor ( id_5416gat, id_5357gat, id_5354gat);
nor ( id_5420gat, id_5301gat, id_5360gat);
nor ( id_5421gat, id_5360gat, id_5298gat);
nor ( id_5422gat, id_5364gat, id_5365gat);
nor ( id_5425gat, id_5309gat, id_5366gat);
nor ( id_5426gat, id_5366gat, id_5241gat);
nor ( id_5427gat, id_5312gat, id_5370gat);
nor ( id_5428gat, id_5370gat, id_5246gat);
nor ( id_5429gat, id_5315gat, id_5374gat);
nor ( id_5430gat, id_5374gat, id_5251gat);
nor ( id_5431gat, id_5378gat, id_5379gat);
nor ( id_5434gat, id_5380gat, id_774gat);
nor ( id_5438gat, id_5324gat, id_5383gat);
nor ( id_5439gat, id_5383gat, id_822gat);
nor ( id_5440gat, id_5200gat, id_5383gat);
nor ( id_5443gat, id_5387gat, id_5388gat);
nor ( id_5446gat, id_5392gat, id_5389gat);
nor ( id_5450gat, id_5336gat, id_5395gat);
nor ( id_5451gat, id_5395gat, id_5333gat);
nor ( id_5452gat, id_5399gat, id_5400gat);
nor ( id_5455gat, id_5401gat, id_1017gat);
nor ( id_5459gat, id_5345gat, id_5404gat);
nor ( id_5460gat, id_5404gat, id_1065gat);
nor ( id_5461gat, id_5221gat, id_5404gat);
nor ( id_5464gat, id_5408gat, id_5409gat);
nor ( id_5467gat, id_5413gat, id_5410gat);
nor ( id_5471gat, id_5357gat, id_5416gat);
nor ( id_5472gat, id_5416gat, id_5354gat);
nor ( id_5473gat, id_5420gat, id_5421gat);
nor ( id_5476gat, id_5422gat, id_1260gat);
nor ( id_5480gat, id_5425gat, id_5426gat);
nor ( id_5483gat, id_5427gat, id_5428gat);
nor ( id_5486gat, id_5429gat, id_5430gat);
nor ( id_5489gat, id_5431gat, id_726gat);
nor ( id_5493gat, id_5380gat, id_5434gat);
nor ( id_5494gat, id_5434gat, id_774gat);
nor ( id_5495gat, id_5262gat, id_5434gat);
nor ( id_5498gat, id_5438gat, id_5439gat);
nor ( id_5501gat, id_5443gat, id_5440gat);
nor ( id_5505gat, id_5392gat, id_5446gat);
nor ( id_5506gat, id_5446gat, id_5389gat);
nor ( id_5507gat, id_5450gat, id_5451gat);
nor ( id_5510gat, id_5452gat, id_969gat);
nor ( id_5514gat, id_5401gat, id_5455gat);
nor ( id_5515gat, id_5455gat, id_1017gat);
nor ( id_5516gat, id_5283gat, id_5455gat);
nor ( id_5519gat, id_5459gat, id_5460gat);
nor ( id_5522gat, id_5464gat, id_5461gat);
nor ( id_5526gat, id_5413gat, id_5467gat);
nor ( id_5527gat, id_5467gat, id_5410gat);
nor ( id_5528gat, id_5471gat, id_5472gat);
nor ( id_5531gat, id_5473gat, id_1212gat);
nor ( id_5535gat, id_5422gat, id_5476gat);
nor ( id_5536gat, id_5476gat, id_1260gat);
nor ( id_5537gat, id_5304gat, id_5476gat);
nor ( id_5540gat, id_5480gat, id_582gat);
nor ( id_5544gat, id_5483gat, id_630gat);
nor ( id_5548gat, id_5486gat, id_678gat);
nor ( id_5552gat, id_5431gat, id_5489gat);
nor ( id_5553gat, id_5489gat, id_726gat);
nor ( id_5554gat, id_5318gat, id_5489gat);
nor ( id_5557gat, id_5493gat, id_5494gat);
nor ( id_5560gat, id_5498gat, id_5495gat);
nor ( id_5564gat, id_5443gat, id_5501gat);
nor ( id_5565gat, id_5501gat, id_5440gat);
nor ( id_5566gat, id_5505gat, id_5506gat);
nor ( id_5569gat, id_5507gat, id_921gat);
nor ( id_5573gat, id_5452gat, id_5510gat);
nor ( id_5574gat, id_5510gat, id_969gat);
nor ( id_5575gat, id_5339gat, id_5510gat);
nor ( id_5578gat, id_5514gat, id_5515gat);
nor ( id_5581gat, id_5519gat, id_5516gat);
nor ( id_5585gat, id_5464gat, id_5522gat);
nor ( id_5586gat, id_5522gat, id_5461gat);
nor ( id_5587gat, id_5526gat, id_5527gat);
nor ( id_5590gat, id_5528gat, id_1164gat);
nor ( id_5594gat, id_5473gat, id_5531gat);
nor ( id_5595gat, id_5531gat, id_1212gat);
nor ( id_5596gat, id_5360gat, id_5531gat);
nor ( id_5599gat, id_5535gat, id_5536gat);
nor ( id_5602gat, id_1308gat, id_5537gat);
nor ( id_5606gat, id_5480gat, id_5540gat);
nor ( id_5607gat, id_5540gat, id_582gat);
nor ( id_5608gat, id_5366gat, id_5540gat);
nor ( id_5611gat, id_5483gat, id_5544gat);
nor ( id_5612gat, id_5544gat, id_630gat);
nor ( id_5613gat, id_5370gat, id_5544gat);
nor ( id_5616gat, id_5486gat, id_5548gat);
nor ( id_5617gat, id_5548gat, id_678gat);
nor ( id_5618gat, id_5374gat, id_5548gat);
nor ( id_5621gat, id_5552gat, id_5553gat);
nor ( id_5624gat, id_5557gat, id_5554gat);
nor ( id_5628gat, id_5498gat, id_5560gat);
nor ( id_5629gat, id_5560gat, id_5495gat);
nor ( id_5630gat, id_5564gat, id_5565gat);
nor ( id_5633gat, id_5566gat, id_873gat);
nor ( id_5637gat, id_5507gat, id_5569gat);
nor ( id_5638gat, id_5569gat, id_921gat);
nor ( id_5639gat, id_5395gat, id_5569gat);
nor ( id_5642gat, id_5573gat, id_5574gat);
nor ( id_5645gat, id_5578gat, id_5575gat);
nor ( id_5649gat, id_5519gat, id_5581gat);
nor ( id_5650gat, id_5581gat, id_5516gat);
nor ( id_5651gat, id_5585gat, id_5586gat);
nor ( id_5654gat, id_5587gat, id_1116gat);
nor ( id_5658gat, id_5528gat, id_5590gat);
nor ( id_5659gat, id_5590gat, id_1164gat);
nor ( id_5660gat, id_5416gat, id_5590gat);
nor ( id_5663gat, id_5594gat, id_5595gat);
nor ( id_5666gat, id_5599gat, id_5596gat);
nor ( id_5670gat, id_1308gat, id_5602gat);
nor ( id_5671gat, id_5602gat, id_5537gat);
nor ( id_5672gat, id_5606gat, id_5607gat);
nor ( id_5673gat, id_5611gat, id_5612gat);
nor ( id_5676gat, id_5616gat, id_5617gat);
nor ( id_5679gat, id_5621gat, id_5618gat);
nor ( id_5683gat, id_5557gat, id_5624gat);
nor ( id_5684gat, id_5624gat, id_5554gat);
nor ( id_5685gat, id_5628gat, id_5629gat);
nor ( id_5688gat, id_5630gat, id_825gat);
nor ( id_5692gat, id_5566gat, id_5633gat);
nor ( id_5693gat, id_5633gat, id_873gat);
nor ( id_5694gat, id_5446gat, id_5633gat);
nor ( id_5697gat, id_5637gat, id_5638gat);
nor ( id_5700gat, id_5642gat, id_5639gat);
nor ( id_5704gat, id_5578gat, id_5645gat);
nor ( id_5705gat, id_5645gat, id_5575gat);
nor ( id_5706gat, id_5649gat, id_5650gat);
nor ( id_5709gat, id_5651gat, id_1068gat);
nor ( id_5713gat, id_5587gat, id_5654gat);
nor ( id_5714gat, id_5654gat, id_1116gat);
nor ( id_5715gat, id_5467gat, id_5654gat);
nor ( id_5718gat, id_5658gat, id_5659gat);
nor ( id_5721gat, id_5663gat, id_5660gat);
nor ( id_5725gat, id_5599gat, id_5666gat);
nor ( id_5726gat, id_5666gat, id_5596gat);
nor ( id_5727gat, id_5670gat, id_5671gat);
nor ( id_5730gat, id_5673gat, id_5608gat);
nor ( id_5734gat, id_5676gat, id_5613gat);
nor ( id_5738gat, id_5621gat, id_5679gat);
nor ( id_5739gat, id_5679gat, id_5618gat);
nor ( id_5740gat, id_5683gat, id_5684gat);
nor ( id_5743gat, id_5685gat, id_777gat);
nor ( id_5747gat, id_5630gat, id_5688gat);
nor ( id_5748gat, id_5688gat, id_825gat);
nor ( id_5749gat, id_5501gat, id_5688gat);
nor ( id_5752gat, id_5692gat, id_5693gat);
nor ( id_5755gat, id_5697gat, id_5694gat);
nor ( id_5759gat, id_5642gat, id_5700gat);
nor ( id_5760gat, id_5700gat, id_5639gat);
nor ( id_5761gat, id_5704gat, id_5705gat);
nor ( id_5764gat, id_5706gat, id_1020gat);
nor ( id_5768gat, id_5651gat, id_5709gat);
nor ( id_5769gat, id_5709gat, id_1068gat);
nor ( id_5770gat, id_5522gat, id_5709gat);
nor ( id_5773gat, id_5713gat, id_5714gat);
nor ( id_5776gat, id_5718gat, id_5715gat);
nor ( id_5780gat, id_5663gat, id_5721gat);
nor ( id_5781gat, id_5721gat, id_5660gat);
nor ( id_5782gat, id_5725gat, id_5726gat);
nor ( id_5785gat, id_5673gat, id_5730gat);
nor ( id_5786gat, id_5730gat, id_5608gat);
nor ( id_5787gat, id_5676gat, id_5734gat);
nor ( id_5788gat, id_5734gat, id_5613gat);
nor ( id_5789gat, id_5738gat, id_5739gat);
nor ( id_5792gat, id_5740gat, id_729gat);
nor ( id_5796gat, id_5685gat, id_5743gat);
nor ( id_5797gat, id_5743gat, id_777gat);
nor ( id_5798gat, id_5560gat, id_5743gat);
nor ( id_5801gat, id_5747gat, id_5748gat);
nor ( id_5804gat, id_5752gat, id_5749gat);
nor ( id_5808gat, id_5697gat, id_5755gat);
nor ( id_5809gat, id_5755gat, id_5694gat);
nor ( id_5810gat, id_5759gat, id_5760gat);
nor ( id_5813gat, id_5761gat, id_972gat);
nor ( id_5817gat, id_5706gat, id_5764gat);
nor ( id_5818gat, id_5764gat, id_1020gat);
nor ( id_5819gat, id_5581gat, id_5764gat);
nor ( id_5822gat, id_5768gat, id_5769gat);
nor ( id_5825gat, id_5773gat, id_5770gat);
nor ( id_5829gat, id_5718gat, id_5776gat);
nor ( id_5830gat, id_5776gat, id_5715gat);
nor ( id_5831gat, id_5780gat, id_5781gat);
nor ( id_5834gat, id_5785gat, id_5786gat);
nor ( id_5837gat, id_5787gat, id_5788gat);
nor ( id_5840gat, id_5789gat, id_681gat);
nor ( id_5844gat, id_5740gat, id_5792gat);
nor ( id_5845gat, id_5792gat, id_729gat);
nor ( id_5846gat, id_5624gat, id_5792gat);
nor ( id_5849gat, id_5796gat, id_5797gat);
nor ( id_5852gat, id_5801gat, id_5798gat);
nor ( id_5856gat, id_5752gat, id_5804gat);
nor ( id_5857gat, id_5804gat, id_5749gat);
nor ( id_5858gat, id_5808gat, id_5809gat);
nor ( id_5861gat, id_5810gat, id_924gat);
nor ( id_5865gat, id_5761gat, id_5813gat);
nor ( id_5866gat, id_5813gat, id_972gat);
nor ( id_5867gat, id_5645gat, id_5813gat);
nor ( id_5870gat, id_5817gat, id_5818gat);
nor ( id_5873gat, id_5822gat, id_5819gat);
nor ( id_5877gat, id_5773gat, id_5825gat);
nor ( id_5878gat, id_5825gat, id_5770gat);
nor ( id_5879gat, id_5829gat, id_5830gat);
nor ( id_5882gat, id_5834gat, id_585gat);
nor ( id_5886gat, id_5837gat, id_633gat);
nor ( id_5890gat, id_5789gat, id_5840gat);
nor ( id_5891gat, id_5840gat, id_681gat);
nor ( id_5892gat, id_5679gat, id_5840gat);
nor ( id_5895gat, id_5844gat, id_5845gat);
nor ( id_5898gat, id_5849gat, id_5846gat);
nor ( id_5902gat, id_5801gat, id_5852gat);
nor ( id_5903gat, id_5852gat, id_5798gat);
nor ( id_5904gat, id_5856gat, id_5857gat);
nor ( id_5907gat, id_5858gat, id_876gat);
nor ( id_5911gat, id_5810gat, id_5861gat);
nor ( id_5912gat, id_5861gat, id_924gat);
nor ( id_5913gat, id_5700gat, id_5861gat);
nor ( id_5916gat, id_5865gat, id_5866gat);
nor ( id_5919gat, id_5870gat, id_5867gat);
nor ( id_5923gat, id_5822gat, id_5873gat);
nor ( id_5924gat, id_5873gat, id_5819gat);
nor ( id_5925gat, id_5877gat, id_5878gat);
nor ( id_5928gat, id_5834gat, id_5882gat);
nor ( id_5929gat, id_5882gat, id_585gat);
nor ( id_5930gat, id_5730gat, id_5882gat);
nor ( id_5933gat, id_5837gat, id_5886gat);
nor ( id_5934gat, id_5886gat, id_633gat);
nor ( id_5935gat, id_5734gat, id_5886gat);
nor ( id_5938gat, id_5890gat, id_5891gat);
nor ( id_5941gat, id_5895gat, id_5892gat);
nor ( id_5945gat, id_5849gat, id_5898gat);
nor ( id_5946gat, id_5898gat, id_5846gat);
nor ( id_5947gat, id_5902gat, id_5903gat);
nor ( id_5950gat, id_5904gat, id_828gat);
nor ( id_5954gat, id_5858gat, id_5907gat);
nor ( id_5955gat, id_5907gat, id_876gat);
nor ( id_5956gat, id_5755gat, id_5907gat);
nor ( id_5959gat, id_5911gat, id_5912gat);
nor ( id_5962gat, id_5916gat, id_5913gat);
nor ( id_5966gat, id_5870gat, id_5919gat);
nor ( id_5967gat, id_5919gat, id_5867gat);
nor ( id_5968gat, id_5923gat, id_5924gat);
nor ( id_5971gat, id_5928gat, id_5929gat);
nor ( id_5972gat, id_5933gat, id_5934gat);
nor ( id_5975gat, id_5938gat, id_5935gat);
nor ( id_5979gat, id_5895gat, id_5941gat);
nor ( id_5980gat, id_5941gat, id_5892gat);
nor ( id_5981gat, id_5945gat, id_5946gat);
nor ( id_5984gat, id_5947gat, id_780gat);
nor ( id_5988gat, id_5904gat, id_5950gat);
nor ( id_5989gat, id_5950gat, id_828gat);
nor ( id_5990gat, id_5804gat, id_5950gat);
nor ( id_5993gat, id_5954gat, id_5955gat);
nor ( id_5996gat, id_5959gat, id_5956gat);
nor ( id_6000gat, id_5916gat, id_5962gat);
nor ( id_6001gat, id_5962gat, id_5913gat);
nor ( id_6002gat, id_5966gat, id_5967gat);
nor ( id_6005gat, id_5972gat, id_5930gat);
nor ( id_6009gat, id_5938gat, id_5975gat);
nor ( id_6010gat, id_5975gat, id_5935gat);
nor ( id_6011gat, id_5979gat, id_5980gat);
nor ( id_6014gat, id_5981gat, id_732gat);
nor ( id_6018gat, id_5947gat, id_5984gat);
nor ( id_6019gat, id_5984gat, id_780gat);
nor ( id_6020gat, id_5852gat, id_5984gat);
nor ( id_6023gat, id_5988gat, id_5989gat);
nor ( id_6026gat, id_5993gat, id_5990gat);
nor ( id_6030gat, id_5959gat, id_5996gat);
nor ( id_6031gat, id_5996gat, id_5956gat);
nor ( id_6032gat, id_6000gat, id_6001gat);
nor ( id_6035gat, id_5972gat, id_6005gat);
nor ( id_6036gat, id_6005gat, id_5930gat);
nor ( id_6037gat, id_6009gat, id_6010gat);
nor ( id_6040gat, id_6011gat, id_684gat);
nor ( id_6044gat, id_5981gat, id_6014gat);
nor ( id_6045gat, id_6014gat, id_732gat);
nor ( id_6046gat, id_5898gat, id_6014gat);
nor ( id_6049gat, id_6018gat, id_6019gat);
nor ( id_6052gat, id_6023gat, id_6020gat);
nor ( id_6056gat, id_5993gat, id_6026gat);
nor ( id_6057gat, id_6026gat, id_5990gat);
nor ( id_6058gat, id_6030gat, id_6031gat);
nor ( id_6061gat, id_6035gat, id_6036gat);
nor ( id_6064gat, id_6037gat, id_636gat);
nor ( id_6068gat, id_6011gat, id_6040gat);
nor ( id_6069gat, id_6040gat, id_684gat);
nor ( id_6070gat, id_5941gat, id_6040gat);
nor ( id_6073gat, id_6044gat, id_6045gat);
nor ( id_6076gat, id_6049gat, id_6046gat);
nor ( id_6080gat, id_6023gat, id_6052gat);
nor ( id_6081gat, id_6052gat, id_6020gat);
nor ( id_6082gat, id_6056gat, id_6057gat);
nor ( id_6085gat, id_6061gat, id_588gat);
nor ( id_6089gat, id_6037gat, id_6064gat);
nor ( id_6090gat, id_6064gat, id_636gat);
nor ( id_6091gat, id_5975gat, id_6064gat);
nor ( id_6094gat, id_6068gat, id_6069gat);
nor ( id_6097gat, id_6073gat, id_6070gat);
nor ( id_6101gat, id_6049gat, id_6076gat);
nor ( id_6102gat, id_6076gat, id_6046gat);
nor ( id_6103gat, id_6080gat, id_6081gat);
nor ( id_6106gat, id_6061gat, id_6085gat);
nor ( id_6107gat, id_6085gat, id_588gat);
nor ( id_6108gat, id_6005gat, id_6085gat);
nor ( id_6111gat, id_6089gat, id_6090gat);
nor ( id_6114gat, id_6094gat, id_6091gat);
nor ( id_6118gat, id_6073gat, id_6097gat);
nor ( id_6119gat, id_6097gat, id_6070gat);
nor ( id_6120gat, id_6101gat, id_6102gat);
nor ( id_6123gat, id_6106gat, id_6107gat);
nor ( id_6124gat, id_6111gat, id_6108gat);
nor ( id_6128gat, id_6094gat, id_6114gat);
nor ( id_6129gat, id_6114gat, id_6091gat);
nor ( id_6130gat, id_6118gat, id_6119gat);
nor ( id_6133gat, id_6111gat, id_6124gat);
nor ( id_6134gat, id_6124gat, id_6108gat);
nor ( id_6135gat, id_6128gat, id_6129gat);
nor ( id_6138gat, id_6133gat, id_6134gat);
not ( id_6141gat, id_6138gat);
not ( id_6146gat, id_6141gat);
nor ( id_6147gat, id_6124gat, id_6141gat);
not ( id_6150gat, id_6146gat);
nor ( id_6151gat, id_6135gat, id_6147gat);
nor ( id_6155gat, id_6135gat, id_6151gat);
nor ( id_6156gat, id_6151gat, id_6147gat);
nor ( id_6157gat, id_6114gat, id_6151gat);
nor ( id_6160gat, id_6155gat, id_6156gat);
nor ( id_6161gat, id_6130gat, id_6157gat);
nor ( id_6165gat, id_6130gat, id_6161gat);
nor ( id_6166gat, id_6161gat, id_6157gat);
nor ( id_6167gat, id_6097gat, id_6161gat);
nor ( id_6170gat, id_6165gat, id_6166gat);
nor ( id_6171gat, id_6120gat, id_6167gat);
nor ( id_6175gat, id_6120gat, id_6171gat);
nor ( id_6176gat, id_6171gat, id_6167gat);
nor ( id_6177gat, id_6076gat, id_6171gat);
nor ( id_6180gat, id_6175gat, id_6176gat);
nor ( id_6181gat, id_6103gat, id_6177gat);
nor ( id_6185gat, id_6103gat, id_6181gat);
nor ( id_6186gat, id_6181gat, id_6177gat);
nor ( id_6187gat, id_6052gat, id_6181gat);
nor ( id_6190gat, id_6185gat, id_6186gat);
nor ( id_6191gat, id_6082gat, id_6187gat);
nor ( id_6195gat, id_6082gat, id_6191gat);
nor ( id_6196gat, id_6191gat, id_6187gat);
nor ( id_6197gat, id_6026gat, id_6191gat);
nor ( id_6200gat, id_6195gat, id_6196gat);
nor ( id_6201gat, id_6058gat, id_6197gat);
nor ( id_6205gat, id_6058gat, id_6201gat);
nor ( id_6206gat, id_6201gat, id_6197gat);
nor ( id_6207gat, id_5996gat, id_6201gat);
nor ( id_6210gat, id_6205gat, id_6206gat);
nor ( id_6211gat, id_6032gat, id_6207gat);
nor ( id_6215gat, id_6032gat, id_6211gat);
nor ( id_6216gat, id_6211gat, id_6207gat);
nor ( id_6217gat, id_5962gat, id_6211gat);
nor ( id_6220gat, id_6215gat, id_6216gat);
nor ( id_6221gat, id_6002gat, id_6217gat);
nor ( id_6225gat, id_6002gat, id_6221gat);
nor ( id_6226gat, id_6221gat, id_6217gat);
nor ( id_6227gat, id_5919gat, id_6221gat);
nor ( id_6230gat, id_6225gat, id_6226gat);
nor ( id_6231gat, id_5968gat, id_6227gat);
nor ( id_6235gat, id_5968gat, id_6231gat);
nor ( id_6236gat, id_6231gat, id_6227gat);
nor ( id_6237gat, id_5873gat, id_6231gat);
nor ( id_6240gat, id_6235gat, id_6236gat);
nor ( id_6241gat, id_5925gat, id_6237gat);
nor ( id_6245gat, id_5925gat, id_6241gat);
nor ( id_6246gat, id_6241gat, id_6237gat);
nor ( id_6247gat, id_5825gat, id_6241gat);
nor ( id_6250gat, id_6245gat, id_6246gat);
nor ( id_6251gat, id_5879gat, id_6247gat);
nor ( id_6255gat, id_5879gat, id_6251gat);
nor ( id_6256gat, id_6251gat, id_6247gat);
nor ( id_6257gat, id_5776gat, id_6251gat);
nor ( id_6260gat, id_6255gat, id_6256gat);
nor ( id_6261gat, id_5831gat, id_6257gat);
nor ( id_6265gat, id_5831gat, id_6261gat);
nor ( id_6266gat, id_6261gat, id_6257gat);
nor ( id_6267gat, id_5721gat, id_6261gat);
nor ( id_6270gat, id_6265gat, id_6266gat);
nor ( id_6271gat, id_5782gat, id_6267gat);
nor ( id_6275gat, id_5782gat, id_6271gat);
nor ( id_6276gat, id_6271gat, id_6267gat);
nor ( id_6277gat, id_5666gat, id_6271gat);
nor ( id_6280gat, id_6275gat, id_6276gat);
nor ( id_6281gat, id_5727gat, id_6277gat);
nor ( id_6285gat, id_5727gat, id_6281gat);
nor ( id_6286gat, id_6281gat, id_6277gat);
nor ( id_6287gat, id_5602gat, id_6281gat);
nor ( id_6288gat, id_6285gat, id_6286gat);

endmodule
