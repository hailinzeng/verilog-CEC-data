module c5315nr
( id_1 ,id_4 ,id_11 ,id_14 ,id_17 ,id_20 ,id_23 ,id_24 ,id_25 ,id_26 ,id_27 ,id_31 ,id_34 ,id_37 ,id_40 ,id_43 ,id_46 ,id_49 ,id_52 ,id_53 ,id_54 ,id_61 ,id_64 ,id_67 ,id_70 ,id_73 ,id_76 ,id_79 ,id_80 ,id_81 ,id_82 ,id_83 ,id_86 ,id_87 ,id_88 ,id_91 ,id_94 ,id_97 ,id_100 ,id_103 ,id_106 ,id_109 ,id_112 ,id_113 ,id_114 ,id_115 ,id_116 ,id_117 ,id_118 ,id_119 ,id_120 ,id_121 ,id_122 ,id_123 ,id_126 ,id_127 ,id_128 ,id_129 ,id_130 ,id_131 ,id_132 ,id_135 ,id_136 ,id_137 ,id_140 ,id_141 ,id_145 ,id_146 ,id_149 ,id_152 ,id_155 ,id_158 ,id_161 ,id_164 ,id_167 ,id_170 ,id_173 ,id_176 ,id_179 ,id_182 ,id_185 ,id_188 ,id_191 ,id_194 ,id_197 ,id_200 ,id_203 ,id_206 ,id_209 ,id_210 ,id_217 ,id_218 ,id_225 ,id_226 ,id_233 ,id_234 ,id_241 ,id_242 ,id_245 ,id_248 ,id_251 ,id_254 ,id_257 ,id_264 ,id_265 ,id_272 ,id_273 ,id_280 ,id_281 ,id_288 ,id_289 ,id_292 ,id_293 ,id_299 ,id_302 ,id_307 ,id_308 ,id_315 ,id_316 ,id_323 ,id_324 ,id_331 ,id_332 ,id_335 ,id_338 ,id_341 ,id_348 ,id_351 ,id_358 ,id_361 ,id_366 ,id_369 ,id_372 ,id_373 ,id_374 ,id_386 ,id_389 ,id_400 ,id_411 ,id_422 ,id_435 ,id_446 ,id_457 ,id_468 ,id_479 ,id_490 ,id_503 ,id_514 ,id_523 ,id_534 ,id_545 ,id_549 ,id_552 ,id_556 ,id_559 ,id_562 ,id_1497 ,id_1689 ,id_1690 ,id_1691 ,id_1694 ,id_2174 ,id_2358 ,id_2824 ,id_3173 ,id_3546 ,id_3548 ,id_3550 ,id_3552 ,id_3717 ,id_3724 ,id_4087 ,id_4088 ,id_4089 ,id_4090 ,id_4091 ,id_4092 ,id_4115 ,id_144 ,id_298 ,id_973 ,id_594 ,id_599 ,id_600 ,id_601 ,id_602 ,id_603 ,id_604 ,id_611 ,id_612 ,id_810 ,id_848 ,id_849 ,id_850 ,id_851 ,id_634 ,id_815 ,id_845 ,id_847 ,id_926 ,id_923 ,id_921 ,id_892 ,id_887 ,id_606 ,id_656 ,id_809 ,id_993 ,id_978 ,id_949 ,id_939 ,id_889 ,id_593 ,id_636 ,id_704 ,id_717 ,id_820 ,id_639 ,id_673 ,id_707 ,id_715 ,id_598 ,id_610 ,id_588 ,id_615 ,id_626 ,id_632 ,id_1002 ,id_1004 ,id_591 ,id_618 ,id_621 ,id_629 ,id_822 ,id_838 ,id_861 ,id_623 ,id_722 ,id_832 ,id_834 ,id_836 ,id_859 ,id_871 ,id_873 ,id_875 ,id_877 ,id_998 ,id_1000 ,id_575 ,id_585 ,id_661 ,id_693 ,id_747 ,id_752 ,id_757 ,id_762 ,id_787 ,id_792 ,id_797 ,id_802 ,id_642 ,id_664 ,id_667 ,id_670 ,id_676 ,id_696 ,id_699 ,id_702 ,id_818 ,id_813 ,id_824 ,id_826 ,id_828 ,id_830 ,id_854 ,id_863 ,id_865 ,id_867 ,id_869 ,id_712 ,id_727 ,id_732 ,id_737 ,id_742 ,id_772 ,id_777 ,id_782 ,id_645 ,id_648 ,id_651 ,id_654 ,id_679 ,id_682 ,id_685 ,id_688 ,id_843 ,id_882 ,id_767 ,id_807 ,id_658 ,id_690  );

input id_1, id_4, id_11, id_14, id_17, id_20, id_23, id_24, id_25, id_26, id_27, id_31, id_34, id_37, id_40, id_43, id_46, id_49, id_52, id_53, id_54, id_61, id_64, id_67, id_70, id_73, id_76, id_79, id_80, id_81, id_82, id_83, id_86, id_87, id_88, id_91, id_94, id_97, id_100, id_103, id_106, id_109, id_112, id_113, id_114, id_115, id_116, id_117, id_118, id_119, id_120, id_121, id_122, id_123, id_126, id_127, id_128, id_129, id_130, id_131, id_132, id_135, id_136, id_137, id_140, id_141, id_145, id_146, id_149, id_152, id_155, id_158, id_161, id_164, id_167, id_170, id_173, id_176, id_179, id_182, id_185, id_188, id_191, id_194, id_197, id_200, id_203, id_206, id_209, id_210, id_217, id_218, id_225, id_226, id_233, id_234, id_241, id_242, id_245, id_248, id_251, id_254, id_257, id_264, id_265, id_272, id_273, id_280, id_281, id_288, id_289, id_292, id_293, id_299, id_302, id_307, id_308, id_315, id_316, id_323, id_324, id_331, id_332, id_335, id_338, id_341, id_348, id_351, id_358, id_361, id_366, id_369, id_372, id_373, id_374, id_386, id_389, id_400, id_411, id_422, id_435, id_446, id_457, id_468, id_479, id_490, id_503, id_514, id_523, id_534, id_545, id_549, id_552, id_556, id_559, id_562, id_1497, id_1689, id_1690, id_1691, id_1694, id_2174, id_2358, id_2824, id_3173, id_3546, id_3548, id_3550, id_3552, id_3717, id_3724, id_4087, id_4088, id_4089, id_4090, id_4091, id_4092, id_4115;

output id_144, id_298, id_973, id_594, id_599, id_600, id_601, id_602, id_603, id_604, id_611, id_612, id_810, id_848, id_849, id_850, id_851, id_634, id_815, id_845, id_847, id_926, id_923, id_921, id_892, id_887, id_606, id_656, id_809, id_993, id_978, id_949, id_939, id_889, id_593, id_636, id_704, id_717, id_820, id_639, id_673, id_707, id_715, id_598, id_610, id_588, id_615, id_626, id_632, id_1002, id_1004, id_591, id_618, id_621, id_629, id_822, id_838, id_861, id_623, id_722, id_832, id_834, id_836, id_859, id_871, id_873, id_875, id_877, id_998, id_1000, id_575, id_585, id_661, id_693, id_747, id_752, id_757, id_762, id_787, id_792, id_797, id_802, id_642, id_664, id_667, id_670, id_676, id_696, id_699, id_702, id_818, id_813, id_824, id_826, id_828, id_830, id_854, id_863, id_865, id_867, id_869, id_712, id_727, id_732, id_737, id_742, id_772, id_777, id_782, id_645, id_648, id_651, id_654, id_679, id_682, id_685, id_688, id_843, id_882, id_767, id_807, id_658, id_690;

buf ( id_144, id_141);
buf ( id_298, id_293);
and ( id_4114, id_135, id_4115);
not ( id_2825, id_2824);
buf ( id_973, id_3173);
not ( id_3547, id_3546);
not ( id_3549, id_3548);
not ( id_3551, id_3550);
not ( id_3553, id_3552);
not ( id_594, id_545);
not ( id_599, id_348);
not ( id_600, id_366);
and ( id_601, id_552, id_562);
not ( id_602, id_549);
not ( id_603, id_545);
not ( id_604, id_545);
not ( id_611, id_338);
not ( id_612, id_358);
nand ( id_633, id_373, id_1);
and ( id_810, id_141, id_145);
not ( id_814, id_3173);
not ( id_816, id_4114);
and ( id_844, id_2825, id_27);
and ( id_846, id_386, id_556);
not ( id_848, id_245);
not ( id_849, id_552);
not ( id_850, id_562);
not ( id_851, id_559);
and ( id_852, id_386, id_559, id_556, id_552);
not ( id_1502, id_1497);
buf ( id_1528, id_1689);
buf ( id_1552, id_1690);
buf ( id_1609, id_1689);
buf ( id_1633, id_1690);
buf ( id_1697, id_137);
buf ( id_1698, id_137);
buf ( id_1701, id_141);
not ( id_2179, id_2174);
buf ( id_2203, id_1691);
buf ( id_2226, id_1694);
buf ( id_2281, id_1691);
buf ( id_2304, id_1694);
buf ( id_2361, id_254);
buf ( id_2370, id_251);
buf ( id_2382, id_251);
buf ( id_2393, id_248);
buf ( id_2405, id_248);
buf ( id_2418, id_4088);
buf ( id_2442, id_4087);
buf ( id_2476, id_4089);
buf ( id_2500, id_4090);
buf ( id_2533, id_210);
buf ( id_2537, id_210);
buf ( id_2541, id_218);
buf ( id_2545, id_218);
buf ( id_2549, id_226);
buf ( id_2553, id_226);
buf ( id_2557, id_234);
buf ( id_2561, id_234);
buf ( id_2627, id_257);
buf ( id_2631, id_257);
buf ( id_2635, id_265);
buf ( id_2639, id_265);
buf ( id_2643, id_273);
buf ( id_2647, id_273);
buf ( id_2651, id_281);
buf ( id_2655, id_281);
buf ( id_2721, id_335);
buf ( id_2734, id_335);
buf ( id_2816, id_206);
and ( id_2822, id_27, id_31);
buf ( id_2826, id_1);
buf ( id_2828, id_2358);
buf ( id_2882, id_293);
buf ( id_2886, id_302);
buf ( id_2890, id_308);
buf ( id_2894, id_308);
buf ( id_2898, id_316);
buf ( id_2902, id_316);
buf ( id_2948, id_324);
buf ( id_2952, id_324);
buf ( id_2956, id_341);
buf ( id_2960, id_341);
buf ( id_2964, id_351);
buf ( id_2968, id_351);
buf ( id_3024, id_257);
buf ( id_3028, id_257);
buf ( id_3032, id_265);
buf ( id_3036, id_265);
buf ( id_3040, id_273);
buf ( id_3044, id_273);
buf ( id_3048, id_281);
buf ( id_3052, id_281);
buf ( id_3092, id_332);
buf ( id_3105, id_332);
buf ( id_3175, id_549);
and ( id_3176, id_31, id_27);
not ( id_3181, id_2358);
buf ( id_3204, id_324);
buf ( id_3208, id_324);
buf ( id_3212, id_341);
buf ( id_3216, id_341);
buf ( id_3220, id_351);
buf ( id_3224, id_351);
buf ( id_3256, id_293);
buf ( id_3260, id_302);
buf ( id_3264, id_308);
buf ( id_3268, id_308);
buf ( id_3272, id_316);
buf ( id_3276, id_316);
buf ( id_3302, id_361);
buf ( id_3314, id_361);
buf ( id_3354, id_210);
buf ( id_3358, id_210);
buf ( id_3362, id_218);
buf ( id_3366, id_218);
buf ( id_3370, id_226);
buf ( id_3374, id_226);
buf ( id_3378, id_234);
buf ( id_3382, id_234);
not ( id_3440, id_324);
buf ( id_3554, id_242);
buf ( id_3555, id_242);
buf ( id_3556, id_254);
buf ( id_3558, id_4088);
buf ( id_3582, id_4087);
buf ( id_3616, id_4092);
buf ( id_3628, id_4091);
buf ( id_3660, id_4089);
buf ( id_3684, id_4090);
not ( id_3721, id_3717);
not ( id_3728, id_3724);
buf ( id_3737, id_4091);
buf ( id_3757, id_4092);
buf ( id_3795, id_4091);
buf ( id_3815, id_4092);
buf ( id_3972, id_4091);
buf ( id_3991, id_4092);
buf ( id_4030, id_4091);
buf ( id_4049, id_4092);
buf ( id_4110, id_299);
buf ( id_4119, id_446);
buf ( id_4127, id_457);
buf ( id_4135, id_468);
buf ( id_4143, id_422);
buf ( id_4151, id_435);
buf ( id_4159, id_389);
buf ( id_4167, id_400);
buf ( id_4175, id_411);
buf ( id_4183, id_374);
buf ( id_4188, id_4);
buf ( id_4276, id_446);
buf ( id_4284, id_457);
buf ( id_4292, id_468);
buf ( id_4300, id_435);
buf ( id_4308, id_389);
buf ( id_4316, id_400);
buf ( id_4324, id_411);
buf ( id_4332, id_422);
buf ( id_4340, id_374);
buf ( id_4631, id_479);
buf ( id_4639, id_490);
buf ( id_4647, id_503);
buf ( id_4655, id_514);
buf ( id_4663, id_523);
buf ( id_4671, id_534);
buf ( id_4676, id_54);
buf ( id_4764, id_479);
buf ( id_4772, id_503);
buf ( id_4780, id_514);
buf ( id_4788, id_523);
buf ( id_4796, id_534);
buf ( id_4804, id_490);
buf ( id_5082, id_361);
buf ( id_5085, id_369);
buf ( id_5090, id_341);
buf ( id_5093, id_351);
buf ( id_5098, id_308);
buf ( id_5101, id_316);
buf ( id_5108, id_293);
buf ( id_5111, id_302);
buf ( id_5332, id_281);
buf ( id_5335, id_289);
buf ( id_5340, id_265);
buf ( id_5343, id_273);
buf ( id_5348, id_234);
buf ( id_5351, id_257);
buf ( id_5356, id_218);
buf ( id_5359, id_226);
buf ( id_5369, id_210);
not ( id_634, id_633);
and ( id_815, id_136, id_814);
not ( id_845, id_844);
not ( id_847, id_846);
buf ( id_926, id_1697);
buf ( id_923, id_1701);
buf ( id_921, id_2826);
and ( id_2979, id_3553, id_514);
or ( id_2999, id_3547, id_514);
buf ( id_892, id_3175);
buf ( id_887, id_4110);
not ( id_606, id_3175);
and ( id_1580, id_170, id_1528, id_1552);
and ( id_1586, id_173, id_1528, id_1552);
and ( id_1592, id_167, id_1528, id_1552);
and ( id_1598, id_164, id_1528, id_1552);
and ( id_1604, id_161, id_1528, id_1552);
nand ( id_656, id_2822, id_140);
and ( id_1668, id_185, id_1609, id_1633);
and ( id_1674, id_158, id_1609, id_1633);
and ( id_1680, id_152, id_1609, id_1633);
and ( id_1686, id_146, id_1609, id_1633);
and ( id_2254, id_170, id_2203, id_2226);
and ( id_2260, id_173, id_2203, id_2226);
and ( id_2266, id_167, id_2203, id_2226);
and ( id_2272, id_164, id_2203, id_2226);
and ( id_2278, id_161, id_2203, id_2226);
and ( id_2339, id_185, id_2281, id_2304);
and ( id_2345, id_158, id_2281, id_2304);
and ( id_2351, id_152, id_2281, id_2304);
and ( id_2357, id_146, id_2281, id_2304);
and ( id_711, id_106, id_3660, id_3684);
and ( id_721, id_61, id_2418, id_2442);
and ( id_726, id_106, id_3558, id_3582);
and ( id_731, id_49, id_3558, id_3582);
and ( id_736, id_103, id_3558, id_3582);
and ( id_741, id_40, id_3558, id_3582);
and ( id_746, id_37, id_3558, id_3582);
and ( id_751, id_20, id_2418, id_2442);
and ( id_756, id_17, id_2418, id_2442);
and ( id_761, id_70, id_2418, id_2442);
and ( id_766, id_64, id_2418, id_2442);
and ( id_771, id_49, id_3660, id_3684);
and ( id_776, id_103, id_3660, id_3684);
and ( id_781, id_40, id_3660, id_3684);
and ( id_786, id_37, id_3660, id_3684);
and ( id_791, id_20, id_2476, id_2500);
and ( id_796, id_17, id_2476, id_2500);
and ( id_801, id_70, id_2476, id_2500);
and ( id_806, id_64, id_2476, id_2500);
not ( id_809, id_2822);
and ( id_3734, id_123, id_3728, id_3717);
and ( id_842, id_3795, id_3815);
and ( id_858, id_61, id_2476, id_2500);
and ( id_881, id_3737, id_3757);
not ( id_4123, id_4119);
not ( id_4131, id_4127);
not ( id_4139, id_4135);
not ( id_4147, id_4143);
not ( id_4155, id_4151);
not ( id_4163, id_4159);
not ( id_4171, id_4167);
not ( id_4179, id_4175);
not ( id_4187, id_4183);
not ( id_4194, id_4188);
not ( id_4282, id_4276);
not ( id_4290, id_4284);
not ( id_4298, id_4292);
not ( id_4306, id_4300);
not ( id_4314, id_4308);
not ( id_4322, id_4316);
not ( id_4330, id_4324);
not ( id_4338, id_4332);
not ( id_4346, id_4340);
buf ( id_1526, id_1697);
not ( id_1540, id_1528);
not ( id_1564, id_1552);
buf ( id_1606, id_1697);
not ( id_1621, id_1609);
not ( id_1645, id_1633);
and ( id_1661, id_179, id_1609, id_1633);
buf ( id_1688, id_2826);
not ( id_4635, id_4631);
not ( id_4643, id_4639);
not ( id_4651, id_4647);
not ( id_4659, id_4655);
not ( id_4667, id_4663);
not ( id_4675, id_4671);
not ( id_4682, id_4676);
not ( id_4770, id_4764);
not ( id_4778, id_4772);
not ( id_4786, id_4780);
not ( id_4794, id_4788);
not ( id_4802, id_4796);
not ( id_4810, id_4804);
buf ( id_2202, id_1698);
not ( id_2215, id_2203);
not ( id_2238, id_2226);
buf ( id_2279, id_1698);
not ( id_2293, id_2281);
not ( id_2316, id_2304);
and ( id_2332, id_179, id_2281, id_2304);
not ( id_2430, id_2418);
not ( id_2454, id_2442);
not ( id_2488, id_2476);
not ( id_2512, id_2500);
not ( id_2536, id_2533);
not ( id_2540, id_2537);
not ( id_2544, id_2541);
not ( id_2548, id_2545);
not ( id_2552, id_2549);
not ( id_2556, id_2553);
not ( id_2560, id_2557);
not ( id_2564, id_2561);
and ( id_2566, id_3553, id_457, id_2537);
and ( id_2572, id_3553, id_468, id_2545);
and ( id_2578, id_3553, id_422, id_2553);
and ( id_2584, id_3553, id_435, id_2561);
and ( id_2590, id_3547, id_2533);
and ( id_2595, id_3547, id_2541);
and ( id_2600, id_3547, id_2549);
and ( id_2605, id_3547, id_2557);
not ( id_2630, id_2627);
not ( id_2634, id_2631);
not ( id_2638, id_2635);
not ( id_2642, id_2639);
not ( id_2646, id_2643);
not ( id_2650, id_2647);
not ( id_2654, id_2651);
not ( id_2658, id_2655);
and ( id_2660, id_3553, id_389, id_2631);
and ( id_2666, id_3553, id_400, id_2639);
and ( id_2672, id_3553, id_411, id_2647);
and ( id_2678, id_3553, id_374, id_2655);
and ( id_2684, id_3547, id_2627);
and ( id_2689, id_3547, id_2635);
and ( id_2694, id_3547, id_2643);
and ( id_2699, id_3547, id_2651);
not ( id_2728, id_2721);
not ( id_2741, id_2734);
and ( id_2748, id_292, id_2721);
and ( id_2750, id_288, id_2721);
and ( id_2752, id_280, id_2721);
and ( id_2754, id_272, id_2721);
and ( id_2756, id_264, id_2721);
and ( id_2758, id_241, id_2734);
and ( id_2760, id_233, id_2734);
and ( id_2762, id_225, id_2734);
and ( id_2764, id_217, id_2734);
and ( id_2766, id_209, id_2734);
buf ( id_2827, id_1701);
not ( id_2838, id_2828);
not ( id_2847, id_2822);
not ( id_2885, id_2882);
not ( id_2889, id_2886);
not ( id_2893, id_2890);
not ( id_2897, id_2894);
not ( id_2901, id_2898);
not ( id_2905, id_2902);
and ( id_2906, id_2393, id_2886);
and ( id_2909, id_2393, id_479, id_2894);
and ( id_2913, id_2393, id_490, id_2902);
and ( id_2918, id_3554, id_2882);
and ( id_2922, id_3554, id_2890);
and ( id_2927, id_3554, id_2898);
not ( id_2951, id_2948);
not ( id_2955, id_2952);
not ( id_2959, id_2956);
not ( id_2963, id_2960);
not ( id_2967, id_2964);
not ( id_2971, id_2968);
and ( id_2973, id_3553, id_503, id_2952);
not ( id_2980, id_2979);
and ( id_2982, id_3553, id_523, id_2960);
and ( id_2988, id_3553, id_534, id_2968);
and ( id_2994, id_3547, id_2948);
and ( id_3001, id_3547, id_2956);
and ( id_3006, id_3547, id_2964);
not ( id_3027, id_3024);
not ( id_3031, id_3028);
not ( id_3035, id_3032);
not ( id_3039, id_3036);
not ( id_3043, id_3040);
not ( id_3047, id_3044);
not ( id_3051, id_3048);
not ( id_3055, id_3052);
and ( id_3056, id_2393, id_389, id_3028);
and ( id_3060, id_2393, id_400, id_3036);
and ( id_3064, id_2393, id_411, id_3044);
and ( id_3068, id_2393, id_374, id_3052);
and ( id_3073, id_3554, id_3024);
and ( id_3078, id_3554, id_3032);
and ( id_3083, id_3554, id_3040);
and ( id_3088, id_3554, id_3048);
not ( id_3099, id_3092);
not ( id_3112, id_3105);
and ( id_3119, id_372, id_3092);
and ( id_3121, id_366, id_3092);
and ( id_3123, id_358, id_3092);
and ( id_3125, id_348, id_3092);
buf ( id_3126, id_338);
and ( id_3128, id_331, id_3105);
and ( id_3130, id_323, id_3105);
and ( id_3132, id_315, id_3105);
and ( id_3134, id_307, id_3105);
and ( id_3136, id_299, id_3105);
not ( id_3187, id_3181);
buf ( id_3193, id_83);
and ( id_3196, id_86, id_3181);
and ( id_3199, id_88, id_3181);
and ( id_3202, id_88, id_3181);
not ( id_3207, id_3204);
not ( id_3211, id_3208);
not ( id_3215, id_3212);
not ( id_3219, id_3216);
not ( id_3223, id_3220);
not ( id_3227, id_3224);
and ( id_3228, id_2405, id_503, id_3208);
and ( id_3232, id_2405, id_514);
and ( id_3234, id_2405, id_523, id_3216);
and ( id_3238, id_2405, id_534, id_3224);
and ( id_3243, id_3555, id_3204);
or ( id_3247, id_3555, id_514);
and ( id_3249, id_3555, id_3212);
and ( id_3253, id_3555, id_3220);
not ( id_3259, id_3256);
not ( id_3263, id_3260);
not ( id_3267, id_3264);
not ( id_3271, id_3268);
not ( id_3275, id_3272);
not ( id_3279, id_3276);
and ( id_3280, id_2405, id_3260);
and ( id_3283, id_2405, id_479, id_3268);
and ( id_3287, id_2405, id_490, id_3276);
and ( id_3292, id_3555, id_3256);
and ( id_3295, id_3555, id_3264);
and ( id_3299, id_3555, id_3272);
not ( id_3305, id_3302);
buf ( id_3306, id_2816);
buf ( id_3310, id_2816);
not ( id_3317, id_3314);
buf ( id_3318, id_2816);
buf ( id_3322, id_2816);
and ( id_3326, id_2405, id_3302);
and ( id_3333, id_2405, id_3314);
not ( id_3357, id_3354);
not ( id_3361, id_3358);
not ( id_3365, id_3362);
not ( id_3369, id_3366);
not ( id_3373, id_3370);
not ( id_3377, id_3374);
not ( id_3381, id_3378);
not ( id_3385, id_3382);
and ( id_3386, id_2393, id_457, id_3358);
and ( id_3390, id_2393, id_468, id_3366);
and ( id_3394, id_2393, id_422, id_3374);
and ( id_3398, id_2393, id_435, id_3382);
and ( id_3403, id_3554, id_3354);
and ( id_3408, id_3554, id_3362);
and ( id_3413, id_3554, id_3370);
and ( id_3418, id_3554, id_3378);
not ( id_5088, id_5082);
not ( id_5089, id_5085);
not ( id_5096, id_5090);
not ( id_5097, id_5093);
buf ( id_3489, id_3440);
buf ( id_3493, id_3440);
not ( id_3570, id_3558);
not ( id_3594, id_3582);
not ( id_3622, id_3616);
not ( id_3632, id_3628);
and ( id_3637, id_97, id_3616);
and ( id_3640, id_94, id_3616);
and ( id_3643, id_97, id_3616);
and ( id_3646, id_94, id_3616);
not ( id_3672, id_3660);
not ( id_3696, id_3684);
not ( id_3745, id_3737);
not ( id_3765, id_3757);
not ( id_3803, id_3795);
not ( id_3823, id_3815);
not ( id_5338, id_5332);
not ( id_5339, id_5335);
not ( id_5346, id_5340);
not ( id_5347, id_5343);
not ( id_5354, id_5348);
not ( id_5355, id_5351);
not ( id_3979, id_3972);
not ( id_3998, id_3991);
not ( id_4037, id_4030);
not ( id_4056, id_4049);
buf ( id_4094, id_4110);
not ( id_5104, id_5098);
not ( id_5105, id_5101);
not ( id_5114, id_5108);
not ( id_5115, id_5111);
not ( id_5362, id_5356);
not ( id_5363, id_5359);
buf ( id_5366, id_2816);
not ( id_5373, id_5369);
buf ( id_993, id_1688);
buf ( id_978, id_1688);
buf ( id_949, id_1688);
buf ( id_939, id_1688);
and ( id_2568, id_457, id_3551, id_2540);
and ( id_2574, id_468, id_3551, id_2548);
and ( id_2580, id_422, id_3551, id_2556);
and ( id_2586, id_435, id_3551, id_2564);
and ( id_2592, id_3549, id_2536);
and ( id_2597, id_3549, id_2544);
and ( id_2602, id_3549, id_2552);
and ( id_2607, id_3549, id_2560);
and ( id_2662, id_389, id_3551, id_2634);
and ( id_2668, id_400, id_3551, id_2642);
and ( id_2674, id_411, id_3551, id_2650);
and ( id_2680, id_374, id_3551, id_2658);
and ( id_2686, id_3549, id_2630);
and ( id_2691, id_3549, id_2638);
and ( id_2696, id_3549, id_2646);
and ( id_2701, id_3549, id_2654);
and ( id_2907, id_2370, id_2889);
and ( id_2910, id_479, id_2370, id_2897);
and ( id_2914, id_490, id_2370, id_2905);
and ( id_2920, id_3556, id_2885);
and ( id_2924, id_3556, id_2893);
and ( id_2929, id_3556, id_2901);
and ( id_2975, id_503, id_3551, id_2955);
and ( id_2984, id_523, id_3551, id_2963);
and ( id_2990, id_534, id_3551, id_2971);
and ( id_2996, id_3549, id_2951);
and ( id_3003, id_3549, id_2959);
and ( id_3008, id_3549, id_2967);
and ( id_3015, id_2980, id_2999);
and ( id_3057, id_389, id_2370, id_3031);
and ( id_3061, id_400, id_2370, id_3039);
and ( id_3065, id_411, id_2370, id_3047);
and ( id_3069, id_374, id_2370, id_3055);
and ( id_3075, id_3556, id_3027);
and ( id_3080, id_3556, id_3035);
and ( id_3085, id_3556, id_3043);
and ( id_3090, id_3556, id_3051);
and ( id_3229, id_503, id_2382, id_3211);
not ( id_3233, id_3232);
and ( id_3235, id_523, id_2382, id_3219);
and ( id_3239, id_534, id_2382, id_3227);
and ( id_3244, id_2361, id_3207);
and ( id_3250, id_2361, id_3215);
and ( id_3254, id_2361, id_3223);
and ( id_3281, id_2382, id_3263);
and ( id_3284, id_479, id_2382, id_3271);
and ( id_3288, id_490, id_2382, id_3279);
and ( id_3293, id_2361, id_3259);
and ( id_3296, id_2361, id_3267);
and ( id_3300, id_2361, id_3275);
and ( id_3327, id_2382, id_3305);
and ( id_3334, id_2382, id_3317);
and ( id_3387, id_457, id_2370, id_3361);
and ( id_3391, id_468, id_2370, id_3369);
and ( id_3395, id_422, id_2370, id_3377);
and ( id_3399, id_435, id_2370, id_3385);
and ( id_3405, id_3556, id_3357);
and ( id_3410, id_3556, id_3365);
and ( id_3415, id_3556, id_3373);
and ( id_3420, id_3556, id_3381);
nand ( id_3422, id_5085, id_5088);
nand ( id_3423, id_5082, id_5089);
nand ( id_3431, id_5093, id_5096);
nand ( id_3432, id_5090, id_5097);
nand ( id_3895, id_5335, id_5338);
nand ( id_3896, id_5332, id_5339);
nand ( id_3904, id_5343, id_5346);
nand ( id_3905, id_5340, id_5347);
nand ( id_3913, id_5351, id_5354);
nand ( id_3914, id_5348, id_5355);
buf ( id_889, id_4094);
nand ( id_5106, id_5101, id_5104);
nand ( id_5107, id_5098, id_5105);
nand ( id_5116, id_5111, id_5114);
nand ( id_5117, id_5108, id_5115);
nand ( id_5364, id_5359, id_5362);
nand ( id_5365, id_5356, id_5363);
not ( id_593, id_4094);
buf ( id_2881, id_2847);
and ( id_1579, id_200, id_1540, id_1552);
and ( id_1585, id_203, id_1540, id_1552);
and ( id_1591, id_197, id_1540, id_1552);
and ( id_1597, id_194, id_1540, id_1552);
and ( id_1603, id_191, id_1540, id_1552);
and ( id_1667, id_182, id_1621, id_1633);
and ( id_1673, id_188, id_1621, id_1633);
and ( id_1679, id_155, id_1621, id_1633);
and ( id_1685, id_149, id_1621, id_1633);
buf ( id_2877, id_2847);
and ( id_2253, id_200, id_2215, id_2226);
and ( id_2259, id_203, id_2215, id_2226);
and ( id_2265, id_197, id_2215, id_2226);
and ( id_2271, id_194, id_2215, id_2226);
and ( id_2277, id_191, id_2215, id_2226);
and ( id_2338, id_182, id_2293, id_2304);
and ( id_2344, id_188, id_2293, id_2304);
and ( id_2350, id_155, id_2293, id_2304);
and ( id_2356, id_149, id_2293, id_2304);
buf ( id_2869, id_2847);
and ( id_710, id_109, id_3672, id_3684);
buf ( id_2873, id_2847);
and ( id_720, id_11, id_2430, id_2442);
and ( id_725, id_109, id_3570, id_3582);
and ( id_730, id_46, id_3570, id_3582);
and ( id_735, id_100, id_3570, id_3582);
and ( id_740, id_91, id_3570, id_3582);
and ( id_745, id_43, id_3570, id_3582);
and ( id_750, id_76, id_2430, id_2442);
and ( id_755, id_73, id_2430, id_2442);
and ( id_760, id_67, id_2430, id_2442);
and ( id_765, id_14, id_2430, id_2442);
and ( id_770, id_46, id_3672, id_3684);
and ( id_775, id_100, id_3672, id_3684);
and ( id_780, id_91, id_3672, id_3684);
and ( id_785, id_43, id_3672, id_3684);
and ( id_790, id_76, id_2488, id_2500);
and ( id_795, id_73, id_2488, id_2500);
and ( id_800, id_67, id_2488, id_2500);
and ( id_805, id_14, id_2488, id_2500);
and ( id_841, id_120, id_3815);
and ( id_857, id_11, id_2488, id_2500);
and ( id_880, id_118, id_3757);
and ( id_1660, id_176, id_1621, id_1633);
and ( id_2331, id_176, id_2293, id_2304);
or ( id_2569, id_2566, id_2568);
or ( id_2575, id_2572, id_2574);
or ( id_2581, id_2578, id_2580);
or ( id_2587, id_2584, id_2586);
or ( id_2593, id_2590, id_2592, id_457);
or ( id_2598, id_2595, id_2597, id_468);
or ( id_2603, id_2600, id_2602, id_422);
or ( id_2608, id_2605, id_2607, id_435);
or ( id_2663, id_2660, id_2662);
or ( id_2669, id_2666, id_2668);
or ( id_2675, id_2672, id_2674);
or ( id_2681, id_2678, id_2680);
or ( id_2687, id_2684, id_2686, id_389);
or ( id_2692, id_2689, id_2691, id_400);
or ( id_2697, id_2694, id_2696, id_411);
or ( id_2702, id_2699, id_2701, id_374);
and ( id_2747, id_289, id_2728);
and ( id_2749, id_281, id_2728);
and ( id_2751, id_273, id_2728);
and ( id_2753, id_265, id_2728);
and ( id_2755, id_257, id_2728);
and ( id_2757, id_234, id_2741);
and ( id_2759, id_226, id_2741);
and ( id_2761, id_218, id_2741);
and ( id_2763, id_210, id_2741);
and ( id_2765, id_206, id_2741);
or ( id_2908, id_2906, id_2907);
or ( id_2911, id_2909, id_2910);
or ( id_2915, id_2913, id_2914);
or ( id_2925, id_2922, id_2924, id_479);
or ( id_2930, id_2927, id_2929, id_490);
or ( id_2933, id_2918, id_2920);
or ( id_2976, id_2973, id_2975);
or ( id_2985, id_2982, id_2984);
or ( id_2991, id_2988, id_2990);
or ( id_2997, id_2994, id_2996, id_503);
or ( id_3004, id_3001, id_3003, id_523);
or ( id_3009, id_3006, id_3008, id_534);
or ( id_3058, id_3056, id_3057);
or ( id_3062, id_3060, id_3061);
or ( id_3066, id_3064, id_3065);
or ( id_3070, id_3068, id_3069);
or ( id_3076, id_3073, id_3075, id_389);
or ( id_3081, id_3078, id_3080, id_400);
or ( id_3086, id_3083, id_3085, id_411);
or ( id_3091, id_3088, id_3090, id_374);
and ( id_3118, id_369, id_3099);
and ( id_3120, id_361, id_3099);
and ( id_3122, id_351, id_3099);
and ( id_3124, id_341, id_3099);
and ( id_3127, id_324, id_3112);
and ( id_3129, id_316, id_3112);
and ( id_3131, id_308, id_3112);
and ( id_3133, id_302, id_3112);
and ( id_3135, id_293, id_3112);
or ( id_3147, id_3099, id_3126);
and ( id_3195, id_87, id_3187);
and ( id_3198, id_34, id_3187);
and ( id_3201, id_34, id_3187);
or ( id_3230, id_3228, id_3229);
or ( id_3236, id_3234, id_3235);
or ( id_3240, id_3238, id_3239);
or ( id_3245, id_3243, id_3244, id_503);
or ( id_3251, id_3249, id_3250, id_523);
or ( id_3255, id_3253, id_3254, id_534);
or ( id_3282, id_3280, id_3281);
or ( id_3285, id_3283, id_3284);
or ( id_3289, id_3287, id_3288);
or ( id_3297, id_3295, id_3296, id_479);
or ( id_3301, id_3299, id_3300, id_490);
not ( id_3309, id_3306);
not ( id_3313, id_3310);
not ( id_3321, id_3318);
not ( id_3325, id_3322);
or ( id_3328, id_3326, id_3327);
and ( id_3329, id_2405, id_446, id_3310);
or ( id_3335, id_3333, id_3334);
and ( id_3336, id_2405, id_446, id_3322);
and ( id_3341, id_3555, id_3306);
and ( id_3345, id_3555, id_3318);
or ( id_3388, id_3386, id_3387);
or ( id_3392, id_3390, id_3391);
or ( id_3396, id_3394, id_3395);
or ( id_3400, id_3398, id_3399);
or ( id_3406, id_3403, id_3405, id_457);
or ( id_3411, id_3408, id_3410, id_468);
or ( id_3416, id_3413, id_3415, id_422);
or ( id_3421, id_3418, id_3420, id_435);
nand ( id_3424, id_3422, id_3423);
nand ( id_3433, id_3431, id_3432);
not ( id_3492, id_3489);
not ( id_3496, id_3493);
and ( id_3780, id_117, id_3745, id_3757);
and ( id_3783, id_126, id_3745, id_3757);
and ( id_3786, id_127, id_3745, id_3757);
and ( id_3789, id_128, id_3745, id_3757);
and ( id_3838, id_131, id_3803, id_3815);
and ( id_3841, id_129, id_3803, id_3815);
and ( id_3844, id_119, id_3803, id_3815);
and ( id_3847, id_130, id_3803, id_3815);
nand ( id_3897, id_3895, id_3896);
nand ( id_3906, id_3904, id_3905);
nand ( id_3915, id_3913, id_3914);
and ( id_4011, id_122, id_3979, id_3991);
and ( id_4014, id_113, id_3979, id_3991);
and ( id_4017, id_53, id_3979, id_3991);
and ( id_4020, id_114, id_3979, id_3991);
and ( id_4023, id_115, id_3979, id_3991);
and ( id_4069, id_52, id_4037, id_4049);
and ( id_4072, id_112, id_4037, id_4049);
and ( id_4075, id_116, id_4037, id_4049);
and ( id_4078, id_121, id_4037, id_4049);
and ( id_4081, id_123, id_4037, id_4049);
nand ( id_5206, id_5116, id_5117);
nand ( id_5209, id_5106, id_5107);
and ( id_5307, id_3233, id_3247);
or ( id_5322, id_3292, id_3293);
not ( id_5372, id_5366);
nand ( id_5375, id_5366, id_5373);
nand ( id_5399, id_5364, id_5365);
not ( id_2813, id_3015);
or ( id_3197, id_3195, id_3196);
or ( id_3200, id_3198, id_3199);
or ( id_3203, id_3201, id_3202);
buf ( id_3194, id_3193);
not ( id_2570, id_2569);
not ( id_2576, id_2575);
not ( id_2582, id_2581);
not ( id_2588, id_2587);
not ( id_2664, id_2663);
not ( id_2670, id_2669);
not ( id_2676, id_2675);
not ( id_2682, id_2681);
or ( id_2767, id_2749, id_2750);
or ( id_2772, id_2751, id_2752);
or ( id_2776, id_2753, id_2754);
or ( id_2780, id_2755, id_2756);
or ( id_2784, id_2757, id_2758);
or ( id_2788, id_2759, id_2760);
or ( id_2794, id_2761, id_2762);
or ( id_2798, id_2763, id_2764);
or ( id_2802, id_2765, id_2766);
not ( id_2912, id_2911);
not ( id_2916, id_2915);
not ( id_2936, id_2908);
not ( id_2977, id_2976);
not ( id_2986, id_2985);
not ( id_2992, id_2991);
not ( id_3059, id_3058);
not ( id_3063, id_3062);
not ( id_3067, id_3066);
not ( id_3071, id_3070);
or ( id_3137, id_3120, id_3121);
or ( id_3139, id_3122, id_3123);
or ( id_3143, id_3124, id_3125);
or ( id_3151, id_3127, id_3128);
or ( id_3155, id_3129, id_3130);
or ( id_3161, id_3131, id_3132);
or ( id_3165, id_3133, id_3134);
or ( id_3167, id_3135, id_3136);
not ( id_3231, id_3230);
not ( id_3237, id_3236);
not ( id_3241, id_3240);
not ( id_3286, id_3285);
not ( id_3290, id_3289);
and ( id_3330, id_446, id_2382, id_3313);
and ( id_3337, id_446, id_2382, id_3325);
and ( id_3342, id_2361, id_3309);
and ( id_3346, id_2361, id_3321);
not ( id_3348, id_3328);
not ( id_3352, id_3335);
not ( id_3389, id_3388);
not ( id_3393, id_3392);
not ( id_3397, id_3396);
not ( id_3401, id_3400);
and ( id_3845, id_3015, id_3803, id_3823);
or ( id_5126, id_3118, id_3119);
or ( id_5178, id_2747, id_2748);
not ( id_5325, id_3282);
nand ( id_5374, id_5369, id_5372);
not ( id_2810, id_2933);
and ( id_635, id_3197, id_3176);
and ( id_2878, id_24, id_2838);
and ( id_2879, id_25, id_2828);
and ( id_2874, id_26, id_2838);
and ( id_2875, id_81, id_2828);
and ( id_703, id_3200, id_3176);
and ( id_2866, id_79, id_2838);
and ( id_2867, id_23, id_2828);
and ( id_2870, id_82, id_2838);
and ( id_2871, id_80, id_2828);
and ( id_716, id_3203, id_3176);
and ( id_819, id_3194, id_3176);
and ( id_1789, id_3147, id_514);
and ( id_2036, id_514, id_3147);
and ( id_2611, id_2570, id_2593);
and ( id_2615, id_2576, id_2598);
and ( id_2619, id_2582, id_2603);
and ( id_2623, id_2588, id_2608);
and ( id_2705, id_2664, id_2687);
and ( id_2709, id_2670, id_2692);
and ( id_2713, id_2676, id_2697);
and ( id_2717, id_2682, id_2702);
and ( id_2939, id_2912, id_2925);
and ( id_2942, id_2916, id_2930);
buf ( id_2945, id_2933);
and ( id_3012, id_2977, id_2997);
and ( id_3018, id_2986, id_3004);
and ( id_3021, id_2992, id_3009);
or ( id_3331, id_3329, id_3330);
or ( id_3338, id_3336, id_3337);
or ( id_3343, id_3341, id_3342, id_446);
or ( id_3347, id_3345, id_3346, id_446);
not ( id_3428, id_3424);
not ( id_3437, id_3433);
and ( id_3514, id_3433, id_3424, id_3489);
and ( id_3836, id_3352, id_3803, id_3823);
and ( id_3852, id_3071, id_3091);
not ( id_5311, id_5307);
not ( id_3901, id_3897);
not ( id_3910, id_3906);
buf ( id_3934, id_3915);
buf ( id_3938, id_3915);
buf ( id_4652, id_3147);
buf ( id_4783, id_3147);
buf ( id_5137, id_3147);
not ( id_5212, id_5206);
not ( id_5213, id_5209);
and ( id_5260, id_3063, id_3081);
and ( id_5263, id_3067, id_3086);
and ( id_5268, id_3401, id_3421);
and ( id_5271, id_3059, id_3076);
and ( id_5276, id_3393, id_3411);
and ( id_5279, id_3397, id_3416);
and ( id_5289, id_3389, id_3406);
and ( id_5296, id_3237, id_3251);
and ( id_5299, id_3241, id_3255);
and ( id_5304, id_3231, id_3245);
and ( id_5312, id_3286, id_3297);
and ( id_5315, id_3290, id_3301);
not ( id_5328, id_5322);
nand ( id_5396, id_5374, id_5375);
not ( id_5403, id_5399);
and ( id_1286, id_446, id_2802);
not ( id_2809, id_2936);
not ( id_597, id_3348);
and ( id_1031, id_2802, id_446);
not ( id_636, id_635);
or ( id_637, id_2878, id_2879, id_2881);
or ( id_671, id_2874, id_2875, id_2877);
not ( id_704, id_703);
or ( id_705, id_2866, id_2867, id_2869);
or ( id_713, id_2870, id_2871, id_2873);
not ( id_717, id_716);
not ( id_820, id_819);
and ( id_1046, id_2798, id_457);
and ( id_1064, id_2794, id_468);
and ( id_1071, id_422, id_2788);
and ( id_1097, id_2784, id_435);
and ( id_1111, id_2780, id_389);
and ( id_1128, id_2776, id_400);
and ( id_1145, id_2772, id_411);
and ( id_1160, id_2767, id_374);
and ( id_1301, id_457, id_2798);
and ( id_1318, id_468, id_2794);
and ( id_1324, id_422, id_2788);
and ( id_1341, id_435, id_2784);
and ( id_1359, id_389, id_2780);
and ( id_1382, id_400, id_2776);
and ( id_1404, id_411, id_2772);
and ( id_1412, id_374, id_2767);
not ( id_1704, id_3167);
not ( id_1712, id_3165);
buf ( id_1724, id_3165);
and ( id_1742, id_3161, id_479);
and ( id_1749, id_490, id_3155);
and ( id_1775, id_3151, id_503);
and ( id_1806, id_3143, id_523);
and ( id_1823, id_3139, id_534);
not ( id_1829, id_3137);
buf ( id_1837, id_3137);
not ( id_1958, id_3167);
not ( id_1966, id_3165);
buf ( id_1978, id_3165);
and ( id_1995, id_479, id_3161);
and ( id_2001, id_490, id_3155);
and ( id_2018, id_503, id_3151);
and ( id_2059, id_523, id_3143);
and ( id_2081, id_534, id_3139);
buf ( id_2089, id_3137);
not ( id_2106, id_3137);
buf ( id_3170, id_3167);
not ( id_3332, id_3331);
not ( id_3339, id_3338);
not ( id_5132, id_5126);
not ( id_5184, id_5178);
not ( id_3853, id_3852);
not ( id_3874, id_3348);
and ( id_4076, id_2936, id_4037, id_4056);
buf ( id_4116, id_2802);
buf ( id_4124, id_2798);
buf ( id_4132, id_2794);
buf ( id_4140, id_2788);
buf ( id_4148, id_2784);
buf ( id_4156, id_2780);
buf ( id_4164, id_2776);
buf ( id_4172, id_2772);
buf ( id_4180, id_2767);
nor ( id_4228, id_422, id_2788);
buf ( id_4279, id_2802);
buf ( id_4287, id_2798);
buf ( id_4295, id_2794);
buf ( id_4303, id_2784);
buf ( id_4311, id_2780);
buf ( id_4319, id_2776);
buf ( id_4327, id_2772);
buf ( id_4335, id_2788);
buf ( id_4343, id_2767);
nor ( id_4348, id_422, id_2788);
nor ( id_4464, id_374, id_2767);
buf ( id_4628, id_3161);
buf ( id_4636, id_3155);
buf ( id_4644, id_3151);
buf ( id_4660, id_3143);
buf ( id_4668, id_3139);
nor ( id_4716, id_490, id_3155);
buf ( id_4767, id_3161);
buf ( id_4775, id_3151);
buf ( id_4791, id_3143);
buf ( id_4799, id_3139);
buf ( id_4807, id_3155);
nor ( id_4812, id_490, id_3155);
buf ( id_5118, id_3139);
buf ( id_5121, id_3143);
buf ( id_5129, id_3137);
buf ( id_5134, id_3151);
buf ( id_5142, id_3161);
buf ( id_5145, id_3155);
buf ( id_5152, id_3167);
buf ( id_5155, id_3165);
buf ( id_5162, id_2788);
buf ( id_5165, id_2784);
buf ( id_5170, id_2798);
buf ( id_5173, id_2794);
buf ( id_5181, id_2802);
buf ( id_5186, id_2772);
buf ( id_5189, id_2767);
buf ( id_5196, id_2780);
buf ( id_5199, id_2776);
nand ( id_5214, id_5209, id_5212);
nand ( id_5215, id_5206, id_5213);
not ( id_5329, id_5325);
nand ( id_5330, id_5325, id_5328);
not ( id_2807, id_2942);
not ( id_2808, id_2939);
not ( id_2811, id_3021);
not ( id_2812, id_3018);
not ( id_2814, id_3012);
not ( id_2626, id_2623);
not ( id_2622, id_2619);
not ( id_2618, id_2615);
not ( id_2614, id_2611);
not ( id_2720, id_2717);
not ( id_2716, id_2713);
not ( id_2712, id_2709);
not ( id_2708, id_2705);
and ( id_639, id_637, id_2827);
and ( id_673, id_671, id_2827);
and ( id_707, id_705, id_2827);
and ( id_715, id_713, id_2827);
and ( id_3731, id_2945, id_3728, id_3721);
not ( id_4658, id_4652);
nand ( id_1777, id_4652, id_4659);
nand ( id_2019, id_4783, id_4786);
not ( id_4787, id_4783);
and ( id_3350, id_3332, id_3343);
and ( id_3353, id_3339, id_3347);
not ( id_5141, id_5137);
and ( id_3513, id_3428, id_3433, id_3492);
and ( id_3516, id_3424, id_3437, id_3496);
and ( id_3517, id_3437, id_3428, id_3493);
and ( id_3778, id_2717, id_3745, id_3765);
and ( id_3781, id_2713, id_3745, id_3765);
and ( id_3784, id_2709, id_3745, id_3765);
and ( id_3787, id_2705, id_3745, id_3765);
and ( id_3839, id_3021, id_3803, id_3823);
and ( id_3842, id_3018, id_3803, id_3823);
not ( id_5266, id_5260);
not ( id_5267, id_5263);
not ( id_5274, id_5268);
not ( id_5275, id_5271);
not ( id_5302, id_5296);
not ( id_5303, id_5299);
not ( id_5310, id_5304);
nand ( id_3891, id_5304, id_5311);
not ( id_3937, id_3934);
not ( id_3941, id_3938);
and ( id_3955, id_3906, id_3897, id_3934);
and ( id_3958, id_3910, id_3901, id_3938);
and ( id_4009, id_2623, id_3979, id_3998);
and ( id_4012, id_2619, id_3979, id_3998);
and ( id_4015, id_2615, id_3979, id_3998);
and ( id_4018, id_2611, id_3979, id_3998);
and ( id_4067, id_3012, id_4037, id_4056);
and ( id_4070, id_2942, id_4037, id_4056);
and ( id_4073, id_2939, id_4037, id_4056);
and ( id_4079, id_2945, id_4037, id_4056);
nand ( id_5239, id_5214, id_5215);
not ( id_5282, id_5276);
not ( id_5283, id_5279);
not ( id_5293, id_5289);
not ( id_5318, id_5312);
not ( id_5319, id_5315);
nand ( id_5331, id_5322, id_5329);
not ( id_5402, id_5396);
nand ( id_5405, id_5396, id_5403);
and ( id_595, id_2807, id_2808, id_2809, id_2810);
and ( id_596, id_2811, id_2812, id_2813, id_2814);
and ( id_607, id_2626, id_2622, id_2618, id_2614);
and ( id_608, id_2720, id_2716, id_2712, id_2708);
buf ( id_1845, id_1724);
buf ( id_1846, id_1742);
buf ( id_2115, id_1978);
buf ( id_2116, id_1995);
not ( id_4122, id_4116);
nand ( id_1022, id_4116, id_4123);
not ( id_4130, id_4124);
nand ( id_1033, id_4124, id_4131);
not ( id_4138, id_4132);
nand ( id_1051, id_4132, id_4139);
not ( id_4146, id_4140);
nand ( id_1079, id_4140, id_4147);
not ( id_4154, id_4148);
nand ( id_1088, id_4148, id_4155);
not ( id_4162, id_4156);
nand ( id_1099, id_4156, id_4163);
not ( id_4170, id_4164);
nand ( id_1115, id_4164, id_4171);
not ( id_4178, id_4172);
nand ( id_1133, id_4172, id_4179);
not ( id_4186, id_4180);
nand ( id_1151, id_4180, id_4187);
not ( id_4234, id_4228);
nand ( id_1276, id_4279, id_4282);
not ( id_4283, id_4279);
nand ( id_1287, id_4287, id_4290);
not ( id_4291, id_4287);
nand ( id_1305, id_4295, id_4298);
not ( id_4299, id_4295);
nand ( id_1330, id_4303, id_4306);
not ( id_4307, id_4303);
nand ( id_1342, id_4311, id_4314);
not ( id_4315, id_4311);
nand ( id_1363, id_4319, id_4322);
not ( id_4323, id_4319);
nand ( id_1388, id_4327, id_4330);
not ( id_4331, id_4327);
nand ( id_1420, id_4335, id_4338);
not ( id_4339, id_4335);
nand ( id_1428, id_4343, id_4346);
not ( id_4347, id_4343);
not ( id_4634, id_4628);
nand ( id_1729, id_4628, id_4635);
not ( id_4642, id_4636);
nand ( id_1757, id_4636, id_4643);
not ( id_4650, id_4644);
nand ( id_1766, id_4644, id_4651);
nand ( id_1776, id_4655, id_4658);
not ( id_4666, id_4660);
nand ( id_1793, id_4660, id_4667);
not ( id_4674, id_4668);
nand ( id_1811, id_4668, id_4675);
buf ( id_1849, id_1742);
buf ( id_1852, id_1742);
buf ( id_1875, id_54);
not ( id_4722, id_4716);
nand ( id_1982, id_4767, id_4770);
not ( id_4771, id_4767);
nand ( id_2007, id_4775, id_4778);
not ( id_4779, id_4775);
nand ( id_2020, id_4780, id_4787);
nand ( id_2040, id_4791, id_4794);
not ( id_4795, id_4791);
nand ( id_2065, id_4799, id_4802);
not ( id_4803, id_4799);
nand ( id_2097, id_4807, id_4810);
not ( id_4811, id_4807);
buf ( id_2119, id_1995);
buf ( id_2122, id_1995);
not ( id_5124, id_5118);
not ( id_5125, id_5121);
nand ( id_3452, id_5129, id_5132);
not ( id_5133, id_5129);
not ( id_5140, id_5134);
nand ( id_3462, id_5134, id_5141);
not ( id_5168, id_5162);
not ( id_5169, id_5165);
not ( id_5176, id_5170);
not ( id_5177, id_5173);
nand ( id_3484, id_5181, id_5184);
not ( id_5185, id_5181);
nor ( id_3515, id_3513, id_3514);
nor ( id_3518, id_3516, id_3517);
not ( id_3857, id_3853);
nand ( id_3860, id_5263, id_5266);
nand ( id_3861, id_5260, id_5267);
nand ( id_3869, id_5271, id_5274);
nand ( id_3870, id_5268, id_5275);
not ( id_3878, id_3874);
nand ( id_3881, id_5299, id_5302);
nand ( id_3882, id_5296, id_5303);
nand ( id_3890, id_5307, id_5310);
and ( id_3954, id_3901, id_3906, id_3937);
and ( id_3957, id_3897, id_3910, id_3941);
and ( id_4021, id_3353, id_3979, id_3998);
not ( id_4099, id_3170);
buf ( id_4236, id_1071);
not ( id_4354, id_4348);
buf ( id_4406, id_1324);
not ( id_4470, id_4464);
buf ( id_4552, id_1412);
buf ( id_4679, id_1829);
buf ( id_4687, id_1704);
buf ( id_4695, id_1704);
buf ( id_4703, id_1712);
buf ( id_4711, id_1712);
buf ( id_4724, id_1749);
not ( id_4818, id_4812);
buf ( id_4855, id_1958);
buf ( id_4865, id_1966);
buf ( id_4870, id_2001);
buf ( id_4913, id_1958);
buf ( id_4923, id_1966);
buf ( id_4951, id_2106);
buf ( id_5006, id_2089);
buf ( id_5039, id_2106);
not ( id_5148, id_5142);
not ( id_5149, id_5145);
not ( id_5158, id_5152);
not ( id_5159, id_5155);
not ( id_5192, id_5186);
not ( id_5193, id_5189);
not ( id_5202, id_5196);
not ( id_5203, id_5199);
nand ( id_5284, id_5279, id_5282);
nand ( id_5285, id_5276, id_5283);
nand ( id_5320, id_5315, id_5318);
nand ( id_5321, id_5312, id_5319);
nand ( id_5386, id_5330, id_5331);
nand ( id_5404, id_5399, id_5402);
and ( id_598, id_595, id_596, id_597);
not ( id_609, id_3350);
nand ( id_1021, id_4119, id_4122);
nand ( id_1032, id_4127, id_4130);
nand ( id_1050, id_4135, id_4138);
nand ( id_1078, id_4143, id_4146);
nand ( id_1087, id_4151, id_4154);
nand ( id_1098, id_4159, id_4162);
nand ( id_1114, id_4167, id_4170);
nand ( id_1132, id_4175, id_4178);
nand ( id_1150, id_4183, id_4186);
nand ( id_1277, id_4276, id_4283);
nand ( id_1288, id_4284, id_4291);
nand ( id_1306, id_4292, id_4299);
nand ( id_1331, id_4300, id_4307);
nand ( id_1343, id_4308, id_4315);
nand ( id_1364, id_4316, id_4323);
nand ( id_1389, id_4324, id_4331);
nand ( id_1421, id_4332, id_4339);
nand ( id_1429, id_4340, id_4347);
nand ( id_1728, id_4631, id_4634);
nand ( id_1756, id_4639, id_4642);
nand ( id_1765, id_4647, id_4650);
nand ( id_1778, id_1776, id_1777);
nand ( id_1792, id_4663, id_4666);
nand ( id_1810, id_4671, id_4674);
nand ( id_1983, id_4764, id_4771);
nand ( id_2008, id_4772, id_4779);
nand ( id_2021, id_2019, id_2020);
nand ( id_2041, id_4788, id_4795);
nand ( id_2066, id_4796, id_4803);
nand ( id_2098, id_4804, id_4811);
nand ( id_3443, id_5121, id_5124);
nand ( id_3444, id_5118, id_5125);
nand ( id_3453, id_5126, id_5133);
nand ( id_3461, id_5137, id_5140);
nand ( id_3466, id_5165, id_5168);
nand ( id_3467, id_5162, id_5169);
nand ( id_3475, id_5173, id_5176);
nand ( id_3476, id_5170, id_5177);
nand ( id_3485, id_5178, id_5185);
not ( id_5243, id_5239);
nand ( id_3862, id_3860, id_3861);
nand ( id_3871, id_3869, id_3870);
nand ( id_3883, id_3881, id_3882);
nand ( id_3892, id_3890, id_3891);
nor ( id_3956, id_3954, id_3955);
nor ( id_3959, id_3957, id_3958);
or ( id_4756, id_1837, id_1875);
nand ( id_5150, id_5145, id_5148);
nand ( id_5151, id_5142, id_5149);
nand ( id_5160, id_5155, id_5158);
nand ( id_5161, id_5152, id_5159);
nand ( id_5194, id_5189, id_5192);
nand ( id_5195, id_5186, id_5193);
nand ( id_5204, id_5199, id_5202);
nand ( id_5205, id_5196, id_5203);
nand ( id_5236, id_3518, id_3515);
buf ( id_5286, id_3350);
nand ( id_5379, id_5284, id_5285);
nand ( id_5389, id_5320, id_5321);
nand ( id_5425, id_5404, id_5405);
and ( id_610, id_607, id_608, id_609);
nand ( id_1023, id_1021, id_1022);
nand ( id_1034, id_1032, id_1033);
nand ( id_1052, id_1050, id_1051);
nand ( id_1080, id_1078, id_1079);
nand ( id_1089, id_1087, id_1088);
nand ( id_1100, id_1098, id_1099);
nand ( id_1116, id_1114, id_1115);
nand ( id_1134, id_1132, id_1133);
nand ( id_1152, id_1150, id_1151);
not ( id_4242, id_4236);
nand ( id_1278, id_1276, id_1277);
nand ( id_1289, id_1287, id_1288);
nand ( id_1307, id_1305, id_1306);
nand ( id_1332, id_1330, id_1331);
nand ( id_1344, id_1342, id_1343);
nand ( id_1365, id_1363, id_1364);
nand ( id_1390, id_1388, id_1389);
nand ( id_1422, id_1420, id_1421);
nand ( id_1430, id_1428, id_1429);
nand ( id_1730, id_1728, id_1729);
nand ( id_1758, id_1756, id_1757);
nand ( id_1767, id_1765, id_1766);
nand ( id_1794, id_1792, id_1793);
nand ( id_1812, id_1810, id_1811);
nand ( id_1876, id_4679, id_4682);
not ( id_4683, id_4679);
not ( id_4691, id_4687);
not ( id_4699, id_4695);
not ( id_4707, id_4703);
not ( id_4715, id_4711);
not ( id_4730, id_4724);
nand ( id_1984, id_1982, id_1983);
nand ( id_2009, id_2007, id_2008);
nand ( id_2042, id_2040, id_2041);
nand ( id_2067, id_2065, id_2066);
nand ( id_2099, id_2097, id_2098);
not ( id_4869, id_4865);
not ( id_4927, id_4923);
nand ( id_3445, id_3443, id_3444);
nand ( id_3454, id_3452, id_3453);
nand ( id_3463, id_3461, id_3462);
nand ( id_3468, id_3466, id_3467);
nand ( id_3477, id_3475, id_3476);
nand ( id_3486, id_3484, id_3485);
not ( id_4412, id_4406);
not ( id_4558, id_4552);
not ( id_4859, id_4855);
not ( id_4876, id_4870);
not ( id_4917, id_4913);
not ( id_4955, id_4951);
not ( id_5012, id_5006);
not ( id_5043, id_5039);
nand ( id_5216, id_5160, id_5161);
nand ( id_5219, id_5150, id_5151);
nand ( id_5226, id_5204, id_5205);
nand ( id_5229, id_5194, id_5195);
not ( id_5392, id_5386);
nand ( id_5422, id_3959, id_3956);
and ( id_1866, id_1778, id_1806);
nand ( id_1877, id_4676, id_4683);
not ( id_4762, id_4756);
and ( id_2142, id_2021, id_2059);
and ( id_2146, id_2021, id_2059);
not ( id_5242, id_5236);
nand ( id_3532, id_5236, id_5243);
not ( id_3866, id_3862);
not ( id_3887, id_3883);
buf ( id_3918, id_3871);
buf ( id_3922, id_3871);
buf ( id_3926, id_3892);
buf ( id_3930, id_3892);
not ( id_5429, id_5425);
buf ( id_4104, id_4099);
buf ( id_4743, id_1778);
buf ( id_4991, id_2021);
buf ( id_5001, id_2021);
not ( id_5292, id_5286);
nand ( id_5295, id_5286, id_5293);
not ( id_5383, id_5379);
not ( id_5393, id_5389);
nand ( id_5394, id_5389, id_5392);
and ( id_1439, id_1278, id_1301);
and ( id_1440, id_1289, id_1278, id_1318);
and ( id_1441, id_1307, id_1278, id_1324, id_1289);
and ( id_1847, id_1730, id_1749);
and ( id_1168, id_1023, id_1046);
and ( id_1169, id_1034, id_1023, id_1064);
and ( id_1170, id_1052, id_1023, id_1071, id_1034);
and ( id_2117, id_1984, id_2001);
not ( id_1086, id_1080);
and ( id_1166, id_1034, id_1080, id_1052, id_1023);
and ( id_1171, id_1034, id_1064);
and ( id_1172, id_1052, id_1071, id_1034);
and ( id_1173, id_1080, id_1052, id_1034);
and ( id_1174, id_1034, id_1064);
and ( id_1175, id_1071, id_1052, id_1034);
and ( id_1176, id_1052, id_1071);
and ( id_1177, id_1080, id_1052);
and ( id_1178, id_1052, id_1071);
and ( id_1179, id_1100, id_1152, id_1116, id_1089, id_1134);
and ( id_1181, id_1089, id_1111);
and ( id_1182, id_1100, id_1089, id_1128);
and ( id_1183, id_1116, id_1089, id_1145, id_1100);
and ( id_1184, id_1134, id_1116, id_1089, id_1160, id_1100);
and ( id_1188, id_1100, id_1128);
and ( id_1189, id_1116, id_1145, id_1100);
and ( id_1190, id_1134, id_1116, id_1160, id_1100);
and ( id_1191, id_4, id_1152, id_1116, id_1134, id_1100);
and ( id_1192, id_1145, id_1116);
and ( id_1193, id_1134, id_1116, id_1160);
and ( id_1194, id_4, id_1152, id_1116, id_1134);
and ( id_1195, id_1134, id_1160);
and ( id_1196, id_4, id_1152, id_1134);
and ( id_1197, id_4, id_1152);
and ( id_1437, id_1422, id_1307, id_1289, id_1278);
and ( id_1442, id_1289, id_1318);
and ( id_1443, id_1307, id_1324, id_1289);
and ( id_1444, id_1422, id_1307, id_1289);
and ( id_1445, id_1289, id_1318);
and ( id_1446, id_1307, id_1324, id_1289);
and ( id_1447, id_1307, id_1324);
and ( id_1451, id_1430, id_1390, id_1365, id_1344, id_1332);
and ( id_1454, id_1332, id_1359);
and ( id_1455, id_1344, id_1332, id_1382);
and ( id_1456, id_1365, id_1332, id_1404, id_1344);
and ( id_1457, id_1390, id_1365, id_1332, id_1412, id_1344);
and ( id_1465, id_1344, id_1382);
and ( id_1466, id_1365, id_1404, id_1344);
and ( id_1467, id_1390, id_1365, id_1412, id_1344);
and ( id_1468, id_1430, id_1365, id_1344, id_1390);
and ( id_1469, id_1344, id_1382);
and ( id_1470, id_1365, id_1404, id_1344);
and ( id_1471, id_1390, id_1365, id_1412, id_1344);
and ( id_1472, id_1365, id_1404);
and ( id_1473, id_1390, id_1365, id_1412);
and ( id_1474, id_1430, id_1365, id_1390);
and ( id_1475, id_1365, id_1404);
and ( id_1476, id_1390, id_1365, id_1412);
and ( id_1477, id_1390, id_1412);
and ( id_1481, id_1422, id_1307);
and ( id_1482, id_1430, id_1390);
not ( id_1764, id_1758);
and ( id_1843, id_1712, id_1758, id_1730, id_1704);
and ( id_1850, id_1730, id_1749);
and ( id_1851, id_1758, id_1730);
and ( id_1853, id_1749, id_1730);
and ( id_1854, id_1730, id_1749);
and ( id_1855, id_1758, id_1730);
and ( id_1856, id_1730, id_1749);
and ( id_1857, id_1778, id_1829, id_1794, id_1767, id_1812);
and ( id_1859, id_1767, id_1789);
and ( id_1860, id_1778, id_1767, id_1806);
and ( id_1861, id_1794, id_1767, id_1823, id_1778);
and ( id_1862, id_1812, id_1794, id_1767, id_1837, id_1778);
and ( id_1867, id_1794, id_1823, id_1778);
and ( id_1868, id_1812, id_1794, id_1837, id_1778);
and ( id_1869, id_54, id_1794, id_1812, id_1778);
and ( id_1870, id_1823, id_1794);
and ( id_1871, id_1812, id_1794, id_1837);
and ( id_1872, id_54, id_1794, id_1812);
and ( id_1873, id_1812, id_1837);
and ( id_1874, id_54, id_1812);
nand ( id_1878, id_1876, id_1877);
and ( id_2113, id_2099, id_1984, id_1966, id_1958);
and ( id_2120, id_1984, id_2001);
and ( id_2121, id_2099, id_1984);
and ( id_2123, id_1984, id_2001);
and ( id_2124, id_1984, id_2001);
and ( id_2128, id_2106, id_2067, id_2042, id_2021, id_2009);
and ( id_2131, id_2009, id_2036);
and ( id_2132, id_2021, id_2009, id_2059);
and ( id_2133, id_2042, id_2009, id_2081, id_2021);
and ( id_2134, id_2067, id_2042, id_2009, id_2089, id_2021);
and ( id_2143, id_2042, id_2081, id_2021);
and ( id_2145, id_2042, id_2021, id_2067);
and ( id_2147, id_2042, id_2081, id_2021);
and ( id_2148, id_2067, id_2042, id_2089, id_2021);
and ( id_2149, id_2042, id_2081);
and ( id_2151, id_2042, id_2067);
and ( id_2152, id_2042, id_2081);
and ( id_2153, id_2067, id_2042, id_2089);
and ( id_2154, id_2067, id_2089);
and ( id_2158, id_2099, id_1984);
buf ( id_2159, id_2067);
not ( id_3449, id_3445);
not ( id_3458, id_3454);
not ( id_3472, id_3468);
not ( id_3481, id_3477);
buf ( id_3497, id_3463);
buf ( id_3501, id_3463);
buf ( id_3505, id_3486);
buf ( id_3509, id_3486);
nand ( id_3531, id_5239, id_5242);
not ( id_5428, id_5422);
nand ( id_3967, id_5422, id_5429);
buf ( id_4191, id_1152);
buf ( id_4199, id_1023);
buf ( id_4207, id_1023);
buf ( id_4215, id_1034);
buf ( id_4223, id_1034);
buf ( id_4231, id_1052);
buf ( id_4239, id_1052);
buf ( id_4247, id_1089);
buf ( id_4255, id_1100);
buf ( id_4263, id_1116);
buf ( id_4271, id_1134);
buf ( id_4371, id_1422);
buf ( id_4381, id_1307);
buf ( id_4391, id_1278);
buf ( id_4401, id_1289);
buf ( id_4429, id_1422);
buf ( id_4439, id_1307);
buf ( id_4449, id_1278);
buf ( id_4459, id_1289);
buf ( id_4497, id_1430);
buf ( id_4507, id_1390);
buf ( id_4517, id_1332);
buf ( id_4527, id_1365);
buf ( id_4537, id_1344);
buf ( id_4547, id_1344);
buf ( id_4585, id_1430);
buf ( id_4595, id_1390);
buf ( id_4605, id_1332);
buf ( id_4615, id_1365);
buf ( id_4719, id_1730);
buf ( id_4727, id_1730);
buf ( id_4735, id_1767);
buf ( id_4751, id_1794);
buf ( id_4759, id_1812);
buf ( id_4835, id_2099);
buf ( id_4845, id_1984);
buf ( id_4893, id_2099);
buf ( id_4903, id_1984);
buf ( id_4961, id_2067);
buf ( id_4971, id_2009);
buf ( id_4981, id_2042);
buf ( id_5049, id_2067);
buf ( id_5059, id_2009);
buf ( id_5069, id_2042);
not ( id_5222, id_5216);
not ( id_5223, id_5219);
not ( id_5232, id_5226);
not ( id_5233, id_5229);
nand ( id_5294, id_5289, id_5292);
nand ( id_5395, id_5386, id_5393);
or ( id_589, id_1286, id_1439, id_1440, id_1441);
or ( id_616, id_3167, id_1845, id_1846, id_1847);
or ( id_619, id_1031, id_1168, id_1169, id_1170);
or ( id_627, id_3167, id_2115, id_2116, id_2117);
or ( id_1185, id_1097, id_1181, id_1182, id_1183, id_1184);
or ( id_1448, id_1318, id_1447);
or ( id_1458, id_1341, id_1454, id_1455, id_1456, id_1457);
or ( id_1478, id_1404, id_1477);
or ( id_1863, id_1775, id_1859, id_1860, id_1861, id_1862);
not ( id_4747, id_4743);
or ( id_2125, id_1995, id_2124);
or ( id_2135, id_2018, id_2131, id_2132, id_2133, id_2134);
or ( id_2155, id_2081, id_2154);
not ( id_4995, id_4991);
not ( id_5005, id_5001);
nand ( id_3533, id_3531, id_3532);
not ( id_3921, id_3918);
not ( id_3925, id_3922);
not ( id_3929, id_3926);
not ( id_3933, id_3930);
and ( id_3943, id_3862, id_3853, id_3918);
and ( id_3946, id_3866, id_3857, id_3922);
and ( id_3949, id_3883, id_3874, id_3926);
and ( id_3952, id_3887, id_3878, id_3930);
nand ( id_3966, id_5425, id_5428);
nand ( id_4107, id_4104, id_132);
or ( id_4196, id_1046, id_1171, id_1172, id_1173);
nor ( id_4204, id_1046, id_1174, id_1175);
or ( id_4212, id_1064, id_1176, id_1177);
nor ( id_4220, id_1064, id_1178);
or ( id_4244, id_1111, id_1188, id_1189, id_1190, id_1191);
or ( id_4252, id_1128, id_1192, id_1193, id_1194);
or ( id_4260, id_1145, id_1195, id_1196);
or ( id_4268, id_1160, id_1197);
or ( id_4361, id_1301, id_1442, id_1443, id_1444);
nor ( id_4419, id_1301, id_1445, id_1446);
or ( id_4467, id_1382, id_1472, id_1473, id_1474);
or ( id_4487, id_1359, id_1465, id_1466, id_1467, id_1468);
nor ( id_4555, id_1382, id_1475, id_1476);
nor ( id_4575, id_1359, id_1469, id_1470, id_1471);
or ( id_4684, id_1724, id_1849, id_1850, id_1851);
nor ( id_4692, id_1724, id_1852, id_1853);
or ( id_4700, id_1742, id_1854, id_1855);
nor ( id_4708, id_1742, id_1856);
or ( id_4732, id_1789, id_1866, id_1867, id_1868, id_1869);
or ( id_4740, id_1806, id_1870, id_1871, id_1872);
or ( id_4748, id_1823, id_1873, id_1874);
or ( id_4825, id_1978, id_2119, id_2120, id_2121);
nor ( id_4883, id_1978, id_2122, id_2123);
or ( id_4928, id_2059, id_2149, id_2151);
or ( id_4941, id_2036, id_2142, id_2143, id_2145);
nor ( id_5009, id_2059, id_2152, id_2153);
nor ( id_5029, id_2036, id_2146, id_2147, id_2148);
nand ( id_5224, id_5219, id_5222);
nand ( id_5225, id_5216, id_5223);
nand ( id_5234, id_5229, id_5232);
nand ( id_5235, id_5226, id_5233);
nand ( id_5376, id_5294, id_5295);
nand ( id_5417, id_5394, id_5395);
not ( id_576, id_1878);
and ( id_588, id_1437, id_1451);
and ( id_615, id_1843, id_1857);
and ( id_626, id_2113, id_2128);
and ( id_632, id_1166, id_1179);
nand ( id_1198, id_4191, id_4194);
not ( id_4195, id_4191);
not ( id_4203, id_4199);
not ( id_4211, id_4207);
not ( id_4219, id_4215);
not ( id_4227, id_4223);
nand ( id_1217, id_4231, id_4234);
not ( id_4235, id_4231);
nand ( id_1221, id_4239, id_4242);
not ( id_4243, id_4239);
and ( id_1224, id_1179, id_4);
not ( id_4251, id_4247);
not ( id_4259, id_4255);
not ( id_4267, id_4263);
not ( id_4275, id_4271);
not ( id_1453, id_1451);
not ( id_4405, id_4401);
not ( id_4463, id_4459);
not ( id_4541, id_4537);
not ( id_4551, id_4547);
nand ( id_1895, id_4719, id_4722);
not ( id_4723, id_4719);
nand ( id_1899, id_4727, id_4730);
not ( id_4731, id_4727);
and ( id_1902, id_1857, id_54);
not ( id_4739, id_4735);
not ( id_4755, id_4751);
nand ( id_1929, id_4759, id_4762);
not ( id_4763, id_4759);
not ( id_2130, id_2128);
not ( id_3500, id_3497);
not ( id_3504, id_3501);
not ( id_3508, id_3505);
not ( id_3512, id_3509);
and ( id_3520, id_3454, id_3445, id_3497);
and ( id_3523, id_3458, id_3449, id_3501);
and ( id_3526, id_3477, id_3468, id_3505);
and ( id_3529, id_3481, id_3472, id_3509);
buf ( id_1002, id_3533);
and ( id_3837, id_1878, id_3795, id_3823);
and ( id_3942, id_3857, id_3862, id_3921);
and ( id_3945, id_3853, id_3866, id_3925);
and ( id_3948, id_3878, id_3883, id_3929);
and ( id_3951, id_3874, id_3887, id_3933);
nand ( id_3968, id_3966, id_3967);
not ( id_4375, id_4371);
not ( id_4385, id_4381);
not ( id_4395, id_4391);
not ( id_4433, id_4429);
not ( id_4443, id_4439);
not ( id_4453, id_4449);
not ( id_4501, id_4497);
not ( id_4511, id_4507);
not ( id_4521, id_4517);
not ( id_4531, id_4527);
not ( id_4619, id_4615);
not ( id_4589, id_4585);
not ( id_4599, id_4595);
not ( id_4609, id_4605);
not ( id_4839, id_4835);
not ( id_4849, id_4845);
not ( id_4897, id_4893);
not ( id_4907, id_4903);
not ( id_4965, id_4961);
not ( id_4975, id_4971);
not ( id_4985, id_4981);
not ( id_5073, id_5069);
not ( id_5053, id_5049);
not ( id_5063, id_5059);
nand ( id_5247, id_5224, id_5225);
nand ( id_5255, id_5234, id_5235);
and ( id_590, id_1437, id_1458);
and ( id_617, id_1863, id_1843);
and ( id_620, id_1185, id_1166);
and ( id_628, id_2113, id_2135);
not ( id_3535, id_3533);
nand ( id_1199, id_4188, id_4195);
not ( id_4202, id_4196);
nand ( id_1204, id_4196, id_4203);
not ( id_4210, id_4204);
nand ( id_1207, id_4204, id_4211);
not ( id_4218, id_4212);
nand ( id_1211, id_4212, id_4219);
not ( id_4226, id_4220);
nand ( id_1214, id_4220, id_4227);
nand ( id_1218, id_4228, id_4235);
nand ( id_1222, id_4236, id_4243);
or ( id_1225, id_1185, id_1224);
not ( id_4250, id_4244);
nand ( id_1237, id_4244, id_4251);
not ( id_4258, id_4252);
nand ( id_1242, id_4252, id_4259);
not ( id_4266, id_4260);
nand ( id_1247, id_4260, id_4267);
not ( id_4274, id_4268);
nand ( id_1252, id_4268, id_4275);
not ( id_1462, id_1458);
not ( id_4690, id_4684);
nand ( id_1882, id_4684, id_4691);
not ( id_4698, id_4692);
nand ( id_1885, id_4692, id_4699);
not ( id_4706, id_4700);
nand ( id_1889, id_4700, id_4707);
not ( id_4714, id_4708);
nand ( id_1892, id_4708, id_4715);
nand ( id_1896, id_4716, id_4723);
nand ( id_1900, id_4724, id_4731);
or ( id_1903, id_1863, id_1902);
not ( id_4738, id_4732);
nand ( id_1915, id_4732, id_4739);
not ( id_4746, id_4740);
nand ( id_1920, id_4740, id_4747);
not ( id_4754, id_4748);
nand ( id_1925, id_4748, id_4755);
nand ( id_1930, id_4756, id_4763);
not ( id_2139, id_2135);
and ( id_3519, id_3449, id_3454, id_3500);
and ( id_3522, id_3445, id_3458, id_3504);
and ( id_3525, id_3472, id_3477, id_3508);
and ( id_3528, id_3468, id_3481, id_3512);
or ( id_3848, id_3836, id_3837, id_3838);
nor ( id_3944, id_3942, id_3943);
nor ( id_3947, id_3945, id_3946);
nor ( id_3950, id_3948, id_3949);
nor ( id_3953, id_3951, id_3952);
not ( id_5421, id_5417);
buf ( id_1004, id_3968);
and ( id_4111, id_4104, id_4107);
and ( id_4112, id_4107, id_132);
or ( id_4351, id_1448, id_1481);
not ( id_4365, id_4361);
not ( id_4409, id_1448);
not ( id_4423, id_4419);
not ( id_4471, id_4467);
nand ( id_4472, id_4467, id_4470);
or ( id_4477, id_1478, id_1482);
not ( id_4491, id_4487);
not ( id_4559, id_4555);
nand ( id_4560, id_4555, id_4558);
not ( id_4565, id_1478);
not ( id_4579, id_4575);
or ( id_4815, id_2125, id_2158);
not ( id_4829, id_4825);
not ( id_4873, id_2125);
not ( id_4887, id_4883);
or ( id_4931, id_2155, id_2159);
not ( id_4934, id_4928);
not ( id_4945, id_4941);
not ( id_5013, id_5009);
nand ( id_5014, id_5009, id_5012);
not ( id_5019, id_2155);
not ( id_5033, id_5029);
not ( id_5382, id_5376);
nand ( id_5385, id_5376, id_5383);
or ( id_591, id_589, id_590);
or ( id_618, id_616, id_617);
or ( id_621, id_619, id_620);
or ( id_629, id_627, id_628);
not ( id_3970, id_3968);
nand ( id_1200, id_1198, id_1199);
nand ( id_1203, id_4199, id_4202);
nand ( id_1206, id_4207, id_4210);
nand ( id_1210, id_4215, id_4218);
nand ( id_1213, id_4223, id_4226);
nand ( id_1219, id_1217, id_1218);
nand ( id_1223, id_1221, id_1222);
nand ( id_1236, id_4247, id_4250);
nand ( id_1241, id_4255, id_4258);
nand ( id_1246, id_4263, id_4266);
nand ( id_1251, id_4271, id_4274);
nand ( id_1881, id_4687, id_4690);
nand ( id_1884, id_4695, id_4698);
nand ( id_1888, id_4703, id_4706);
nand ( id_1891, id_4711, id_4714);
nand ( id_1897, id_1895, id_1896);
nand ( id_1901, id_1899, id_1900);
nand ( id_1914, id_4735, id_4738);
nand ( id_1919, id_4743, id_4746);
nand ( id_1924, id_4751, id_4754);
nand ( id_1931, id_1929, id_1930);
nor ( id_3521, id_3519, id_3520);
nor ( id_3524, id_3522, id_3523);
nor ( id_3527, id_3525, id_3526);
nor ( id_3530, id_3528, id_3529);
not ( id_5251, id_5247);
not ( id_5259, id_5255);
or ( id_4113, id_4111, id_4112);
nand ( id_4473, id_4464, id_4471);
nand ( id_4561, id_4552, id_4559);
nand ( id_5015, id_5006, id_5013);
nand ( id_5384, id_5379, id_5382);
nand ( id_5406, id_3947, id_3944);
nand ( id_5414, id_3953, id_3950);
and ( id_1664, id_3848, id_1621, id_1645);
and ( id_2335, id_3848, id_2293, id_2316);
and ( id_718, id_3848, id_2430, id_2454);
not ( id_822, id_3848);
and ( id_855, id_3848, id_2488, id_2512);
nand ( id_1205, id_1203, id_1204);
nand ( id_1208, id_1206, id_1207);
nand ( id_1212, id_1210, id_1211);
nand ( id_1215, id_1213, id_1214);
not ( id_1220, id_1219);
not ( id_1231, id_1225);
nand ( id_1238, id_1236, id_1237);
nand ( id_1243, id_1241, id_1242);
nand ( id_1248, id_1246, id_1247);
nand ( id_1253, id_1251, id_1252);
and ( id_1272, id_1225, id_1086);
and ( id_1483, id_1462, id_1453);
nand ( id_1883, id_1881, id_1882);
nand ( id_1886, id_1884, id_1885);
nand ( id_1890, id_1888, id_1889);
nand ( id_1893, id_1891, id_1892);
not ( id_1898, id_1897);
not ( id_1909, id_1903);
nand ( id_1916, id_1914, id_1915);
nand ( id_1921, id_1919, id_1920);
nand ( id_1926, id_1924, id_1925);
and ( id_1953, id_1903, id_1764);
and ( id_2160, id_2139, id_2130);
not ( id_4355, id_4351);
nand ( id_4356, id_4351, id_4354);
not ( id_4413, id_4409);
nand ( id_4414, id_4409, id_4412);
nand ( id_4474, id_4472, id_4473);
not ( id_4481, id_4477);
nand ( id_4562, id_4560, id_4561);
not ( id_4569, id_4565);
not ( id_4819, id_4815);
nand ( id_4820, id_4815, id_4818);
not ( id_4877, id_4873);
nand ( id_4878, id_4873, id_4876);
not ( id_4935, id_4931);
nand ( id_4936, id_4931, id_4934);
nand ( id_5016, id_5014, id_5015);
not ( id_5023, id_5019);
nand ( id_5244, id_3524, id_3521);
nand ( id_5252, id_3530, id_3527);
nand ( id_5409, id_5384, id_5385);
not ( id_566, id_1200);
not ( id_577, id_1931);
and ( id_3733, id_4113, id_3724, id_3721);
not ( id_1209, id_1208);
not ( id_1216, id_1215);
and ( id_1257, id_1225, id_1205);
and ( id_1262, id_1225, id_1212);
and ( id_1267, id_1225, id_1220);
not ( id_1887, id_1886);
not ( id_1894, id_1893);
and ( id_1935, id_1903, id_1883);
and ( id_1943, id_1903, id_1890);
and ( id_1948, id_1903, id_1898);
and ( id_3779, id_1200, id_3737, id_3765);
and ( id_3840, id_1931, id_3795, id_3823);
not ( id_5412, id_5406);
not ( id_5420, id_5414);
nand ( id_3964, id_5414, id_5421);
nand ( id_4357, id_4348, id_4355);
nand ( id_4415, id_4406, id_4413);
nand ( id_4821, id_4812, id_4819);
nand ( id_4879, id_4870, id_4877);
nand ( id_4937, id_4928, id_4935);
not ( id_567, id_1253);
not ( id_568, id_1248);
not ( id_569, id_1243);
not ( id_570, id_1238);
not ( id_578, id_1926);
not ( id_579, id_1921);
not ( id_580, id_1916);
and ( id_1256, id_1209, id_1231);
and ( id_1261, id_1216, id_1231);
and ( id_1266, id_1223, id_1231);
and ( id_1271, id_1080, id_1231);
not ( id_1486, id_1483);
and ( id_1934, id_1887, id_1909);
and ( id_1942, id_1894, id_1909);
and ( id_1947, id_1901, id_1909);
and ( id_1952, id_1758, id_1909);
not ( id_2163, id_2160);
not ( id_5250, id_5244);
nand ( id_3537, id_5244, id_5251);
not ( id_5258, id_5252);
nand ( id_3542, id_5252, id_5259);
and ( id_3782, id_1253, id_3737, id_3765);
and ( id_3785, id_1248, id_3737, id_3765);
and ( id_3788, id_1243, id_3737, id_3765);
or ( id_3790, id_3778, id_3779, id_3780);
and ( id_3843, id_1926, id_3795, id_3823);
and ( id_3846, id_1921, id_3795, id_3823);
or ( id_3849, id_3839, id_3840, id_3841);
nand ( id_3960, id_5409, id_5412);
not ( id_5413, id_5409);
nand ( id_3963, id_5417, id_5420);
and ( id_4010, id_1238, id_3972, id_3998);
and ( id_4068, id_1916, id_4030, id_4056);
nand ( id_4358, id_4356, id_4357);
nand ( id_4416, id_4414, id_4415);
not ( id_4480, id_4474);
nand ( id_4483, id_4474, id_4481);
not ( id_4568, id_4562);
nand ( id_4571, id_4562, id_4569);
nand ( id_4822, id_4820, id_4821);
nand ( id_4880, id_4878, id_4879);
nand ( id_4938, id_4936, id_4937);
not ( id_5022, id_5016);
nand ( id_5025, id_5016, id_5023);
or ( id_1258, id_1256, id_1257);
or ( id_1263, id_1261, id_1262);
or ( id_1268, id_1266, id_1267);
or ( id_1273, id_1271, id_1272);
or ( id_1936, id_1934, id_1935);
or ( id_1944, id_1942, id_1943);
or ( id_1949, id_1947, id_1948);
or ( id_1954, id_1952, id_1953);
nand ( id_3536, id_5247, id_5250);
nand ( id_3541, id_5255, id_5258);
or ( id_3791, id_3781, id_3782, id_3783);
or ( id_3792, id_3784, id_3785, id_3786);
or ( id_3793, id_3787, id_3788, id_3789);
or ( id_3850, id_3842, id_3843, id_3844);
or ( id_3851, id_3845, id_3846, id_3847);
nand ( id_3961, id_5406, id_5413);
nand ( id_3965, id_3963, id_3964);
or ( id_4024, id_4009, id_4010, id_4011);
or ( id_4082, id_4067, id_4068, id_4069);
nand ( id_4482, id_4477, id_4480);
nand ( id_4570, id_4565, id_4568);
nand ( id_5024, id_5019, id_5022);
and ( id_1666, id_3790, id_1609, id_1645);
and ( id_1670, id_3849, id_1621, id_1645);
and ( id_2337, id_3790, id_2281, id_2316);
and ( id_2341, id_3849, id_2293, id_2316);
and ( id_719, id_3790, id_2418, id_2454);
and ( id_758, id_3849, id_2430, id_2454);
and ( id_798, id_3849, id_2488, id_2512);
not ( id_838, id_3849);
and ( id_856, id_3790, id_2476, id_2512);
not ( id_861, id_3790);
nand ( id_3538, id_3536, id_3537);
nand ( id_3543, id_3541, id_3542);
nand ( id_3962, id_3960, id_3961);
not ( id_4364, id_4358);
nand ( id_4367, id_4358, id_4365);
not ( id_4422, id_4416);
nand ( id_4425, id_4416, id_4423);
nand ( id_4484, id_4482, id_4483);
nand ( id_4572, id_4570, id_4571);
not ( id_4828, id_4822);
nand ( id_4831, id_4822, id_4829);
not ( id_4886, id_4880);
nand ( id_4889, id_4880, id_4887);
not ( id_4944, id_4938);
nand ( id_4947, id_4938, id_4945);
nand ( id_5026, id_5024, id_5025);
not ( id_571, id_1273);
not ( id_572, id_1268);
not ( id_573, id_1263);
not ( id_574, id_1258);
not ( id_581, id_1954);
not ( id_582, id_1949);
not ( id_583, id_1944);
not ( id_584, id_1936);
not ( id_623, id_1936);
and ( id_1576, id_4082, id_1540, id_1564);
and ( id_1578, id_4024, id_1528, id_1564);
or ( id_659, id_1664, id_1666, id_1667, id_1668);
and ( id_1672, id_3791, id_1609, id_1645);
and ( id_1676, id_3850, id_1621, id_1645);
and ( id_1678, id_3792, id_1609, id_1645);
and ( id_1682, id_3851, id_1621, id_1645);
and ( id_1684, id_3793, id_1609, id_1645);
and ( id_2250, id_4082, id_2215, id_2238);
and ( id_2252, id_4024, id_2203, id_2238);
or ( id_691, id_2335, id_2337, id_2338, id_2339);
and ( id_2343, id_3791, id_2281, id_2316);
and ( id_2347, id_3850, id_2293, id_2316);
and ( id_2349, id_3792, id_2281, id_2316);
and ( id_2353, id_3851, id_2293, id_2316);
and ( id_2355, id_3793, id_2281, id_2316);
or ( id_722, id_718, id_719, id_720, id_721);
and ( id_743, id_4082, id_3570, id_3594);
and ( id_744, id_4024, id_3558, id_3594);
and ( id_748, id_3851, id_2430, id_2454);
and ( id_749, id_3793, id_2418, id_2454);
and ( id_753, id_3850, id_2430, id_2454);
and ( id_754, id_3792, id_2418, id_2454);
and ( id_759, id_3791, id_2418, id_2454);
and ( id_783, id_4082, id_3672, id_3696);
and ( id_784, id_4024, id_3660, id_3696);
and ( id_788, id_3851, id_2488, id_2512);
and ( id_789, id_3793, id_2476, id_2512);
and ( id_793, id_3850, id_2488, id_2512);
and ( id_794, id_3792, id_2476, id_2512);
and ( id_799, id_3791, id_2476, id_2512);
and ( id_3735, id_1936, id_3724, id_3717);
not ( id_832, id_4082);
not ( id_834, id_3851);
not ( id_836, id_3850);
not ( id_3835, id_3965);
or ( id_859, id_855, id_856, id_857, id_858);
not ( id_871, id_4024);
not ( id_873, id_3793);
not ( id_875, id_3792);
not ( id_877, id_3791);
buf ( id_998, id_3538);
buf ( id_1000, id_3543);
and ( id_3651, id_3965, id_3632);
and ( id_4013, id_1273, id_3972, id_3998);
and ( id_4016, id_1268, id_3972, id_3998);
and ( id_4019, id_1263, id_3972, id_3998);
and ( id_4022, id_1258, id_3972, id_3998);
and ( id_4071, id_1954, id_4030, id_4056);
and ( id_4074, id_1949, id_4030, id_4056);
and ( id_4077, id_1944, id_4030, id_4056);
and ( id_4080, id_1936, id_4030, id_4056);
nand ( id_4096, id_4113, id_1936);
nand ( id_4366, id_4361, id_4364);
nand ( id_4424, id_4419, id_4422);
nand ( id_4830, id_4825, id_4828);
nand ( id_4888, id_4883, id_4886);
nand ( id_4946, id_4941, id_4944);
and ( id_575, id_566, id_567, id_568, id_569, id_570, id_571, id_572, id_573, id_574);
and ( id_585, id_576, id_577, id_578, id_579, id_580, id_581, id_582, id_583, id_584);
or ( id_640, id_1576, id_1578, id_1579, id_1580);
and ( id_661, id_659, id_1606);
or ( id_662, id_1670, id_1672, id_1673, id_1674);
or ( id_665, id_1676, id_1678, id_1679, id_1680);
or ( id_668, id_1682, id_1684, id_1685, id_1686);
or ( id_674, id_2250, id_2252, id_2253, id_2254);
and ( id_693, id_691, id_2279);
or ( id_694, id_2341, id_2343, id_2344, id_2345);
or ( id_697, id_2347, id_2349, id_2350, id_2351);
or ( id_700, id_2353, id_2355, id_2356, id_2357);
or ( id_747, id_743, id_744, id_745, id_746);
or ( id_752, id_748, id_749, id_750, id_751);
or ( id_757, id_753, id_754, id_755, id_756);
or ( id_762, id_758, id_759, id_760, id_761);
or ( id_787, id_783, id_784, id_785, id_786);
or ( id_792, id_788, id_789, id_790, id_791);
or ( id_797, id_793, id_794, id_795, id_796);
or ( id_802, id_798, id_799, id_800, id_801);
or ( id_817, id_3731, id_3733, id_3734, id_3735);
and ( id_839, id_3835, id_3803, id_3823);
not ( id_3540, id_3538);
not ( id_3545, id_3543);
not ( id_3777, id_3962);
and ( id_3648, id_3962, id_3632);
or ( id_4025, id_4012, id_4013, id_4014);
or ( id_4026, id_4015, id_4016, id_4017);
or ( id_4027, id_4018, id_4019, id_4020);
or ( id_4028, id_4021, id_4022, id_4023);
or ( id_4083, id_4070, id_4071, id_4072);
or ( id_4084, id_4073, id_4074, id_4075);
or ( id_4085, id_4076, id_4077, id_4078);
or ( id_4086, id_4079, id_4080, id_4081);
nand ( id_4368, id_4366, id_4367);
nand ( id_4426, id_4424, id_4425);
not ( id_4490, id_4484);
nand ( id_4493, id_4484, id_4491);
not ( id_4578, id_4572);
nand ( id_4581, id_4572, id_4579);
nand ( id_4832, id_4830, id_4831);
nand ( id_4890, id_4888, id_4889);
nand ( id_4948, id_4946, id_4947);
not ( id_5032, id_5026);
nand ( id_5035, id_5026, id_5033);
and ( id_642, id_640, id_1526);
and ( id_664, id_662, id_1606);
and ( id_667, id_665, id_1606);
and ( id_670, id_668, id_1606);
and ( id_676, id_674, id_2202);
and ( id_696, id_694, id_2279);
and ( id_699, id_697, id_2279);
and ( id_702, id_700, id_2279);
and ( id_811, id_4113, id_4096);
and ( id_812, id_4096, id_1936);
and ( id_818, id_816, id_817);
and ( id_853, id_562, id_3540, id_3545, id_3535, id_3970);
and ( id_878, id_3777, id_3745, id_3765);
nand ( id_4492, id_4487, id_4490);
nand ( id_4580, id_4575, id_4578);
nand ( id_5034, id_5029, id_5032);
and ( id_1582, id_4083, id_1540, id_1564);
and ( id_1584, id_4025, id_1528, id_1564);
and ( id_1588, id_4084, id_1540, id_1564);
and ( id_1590, id_4026, id_1528, id_1564);
and ( id_1594, id_4085, id_1540, id_1564);
and ( id_1596, id_4027, id_1528, id_1564);
and ( id_1600, id_4086, id_1540, id_1564);
and ( id_1602, id_4028, id_1528, id_1564);
and ( id_2256, id_4083, id_2215, id_2238);
and ( id_2258, id_4025, id_2203, id_2238);
and ( id_2262, id_4084, id_2215, id_2238);
and ( id_2264, id_4026, id_2203, id_2238);
and ( id_2268, id_4085, id_2215, id_2238);
and ( id_2270, id_4027, id_2203, id_2238);
and ( id_2274, id_4086, id_2215, id_2238);
and ( id_2276, id_4028, id_2203, id_2238);
and ( id_708, id_4086, id_3672, id_3696);
and ( id_709, id_4028, id_3660, id_3696);
and ( id_723, id_4086, id_3570, id_3594);
and ( id_724, id_4028, id_3558, id_3594);
and ( id_728, id_4085, id_3570, id_3594);
and ( id_729, id_4027, id_3558, id_3594);
and ( id_733, id_4084, id_3570, id_3594);
and ( id_734, id_4026, id_3558, id_3594);
and ( id_738, id_4083, id_3570, id_3594);
and ( id_739, id_4025, id_3558, id_3594);
and ( id_768, id_4085, id_3672, id_3696);
and ( id_769, id_4027, id_3660, id_3696);
and ( id_773, id_4084, id_3672, id_3696);
and ( id_774, id_4026, id_3660, id_3696);
and ( id_778, id_4083, id_3672, id_3696);
and ( id_779, id_4025, id_3660, id_3696);
or ( id_813, id_811, id_812);
not ( id_824, id_4086);
not ( id_826, id_4085);
not ( id_828, id_4084);
not ( id_830, id_4083);
and ( id_854, id_852, id_853, id_245);
not ( id_863, id_4028);
not ( id_865, id_4027);
not ( id_867, id_4026);
not ( id_869, id_4025);
not ( id_4374, id_4368);
nand ( id_4377, id_4368, id_4375);
not ( id_4432, id_4426);
nand ( id_4435, id_4426, id_4433);
nand ( id_4494, id_4492, id_4493);
nand ( id_4582, id_4580, id_4581);
not ( id_4838, id_4832);
nand ( id_4841, id_4832, id_4839);
not ( id_4896, id_4890);
nand ( id_4899, id_4890, id_4897);
not ( id_4954, id_4948);
nand ( id_4957, id_4948, id_4955);
nand ( id_5036, id_5034, id_5035);
or ( id_643, id_1582, id_1584, id_1585, id_1586);
or ( id_646, id_1588, id_1590, id_1591, id_1592);
or ( id_649, id_1594, id_1596, id_1597, id_1598);
or ( id_652, id_1600, id_1602, id_1603, id_1604);
or ( id_677, id_2256, id_2258, id_2259, id_2260);
or ( id_680, id_2262, id_2264, id_2265, id_2266);
or ( id_683, id_2268, id_2270, id_2271, id_2272);
or ( id_686, id_2274, id_2276, id_2277, id_2278);
or ( id_712, id_708, id_709, id_710, id_711);
or ( id_727, id_723, id_724, id_725, id_726);
or ( id_732, id_728, id_729, id_730, id_731);
or ( id_737, id_733, id_734, id_735, id_736);
or ( id_742, id_738, id_739, id_740, id_741);
or ( id_772, id_768, id_769, id_770, id_771);
or ( id_777, id_773, id_774, id_775, id_776);
or ( id_782, id_778, id_779, id_780, id_781);
nand ( id_4376, id_4371, id_4374);
nand ( id_4434, id_4429, id_4432);
nand ( id_4840, id_4835, id_4838);
nand ( id_4898, id_4893, id_4896);
nand ( id_4956, id_4951, id_4954);
and ( id_645, id_643, id_1526);
and ( id_648, id_646, id_1526);
and ( id_651, id_649, id_1526);
and ( id_654, id_652, id_1526);
and ( id_679, id_677, id_2202);
and ( id_682, id_680, id_2202);
and ( id_685, id_683, id_2202);
and ( id_688, id_686, id_2202);
nand ( id_4378, id_4376, id_4377);
nand ( id_4436, id_4434, id_4435);
not ( id_4500, id_4494);
nand ( id_4503, id_4494, id_4501);
not ( id_4588, id_4582);
nand ( id_4591, id_4582, id_4589);
nand ( id_4842, id_4840, id_4841);
nand ( id_4900, id_4898, id_4899);
nand ( id_4958, id_4956, id_4957);
not ( id_5042, id_5036);
nand ( id_5045, id_5036, id_5043);
nand ( id_4502, id_4497, id_4500);
nand ( id_4590, id_4585, id_4588);
nand ( id_5044, id_5039, id_5042);
not ( id_4384, id_4378);
nand ( id_4387, id_4378, id_4385);
not ( id_4442, id_4436);
nand ( id_4445, id_4436, id_4443);
nand ( id_4504, id_4502, id_4503);
nand ( id_4592, id_4590, id_4591);
not ( id_4848, id_4842);
nand ( id_4851, id_4842, id_4849);
not ( id_4906, id_4900);
nand ( id_4909, id_4900, id_4907);
not ( id_4964, id_4958);
nand ( id_4967, id_4958, id_4965);
nand ( id_5046, id_5044, id_5045);
nand ( id_4386, id_4381, id_4384);
nand ( id_4444, id_4439, id_4442);
nand ( id_4850, id_4845, id_4848);
nand ( id_4908, id_4903, id_4906);
nand ( id_4966, id_4961, id_4964);
nand ( id_4388, id_4386, id_4387);
nand ( id_4446, id_4444, id_4445);
not ( id_4510, id_4504);
nand ( id_4513, id_4504, id_4511);
not ( id_4598, id_4592);
nand ( id_4601, id_4592, id_4599);
nand ( id_4852, id_4850, id_4851);
nand ( id_4910, id_4908, id_4909);
nand ( id_4968, id_4966, id_4967);
not ( id_5052, id_5046);
nand ( id_5055, id_5046, id_5053);
nand ( id_4512, id_4507, id_4510);
nand ( id_4600, id_4595, id_4598);
nand ( id_5054, id_5049, id_5052);
not ( id_4394, id_4388);
nand ( id_4397, id_4388, id_4395);
not ( id_4452, id_4446);
nand ( id_4455, id_4446, id_4453);
nand ( id_4514, id_4512, id_4513);
nand ( id_4602, id_4600, id_4601);
not ( id_4858, id_4852);
nand ( id_4861, id_4852, id_4859);
not ( id_4916, id_4910);
nand ( id_4919, id_4910, id_4917);
not ( id_4974, id_4968);
nand ( id_4977, id_4968, id_4975);
nand ( id_5056, id_5054, id_5055);
nand ( id_4396, id_4391, id_4394);
nand ( id_4454, id_4449, id_4452);
nand ( id_4860, id_4855, id_4858);
nand ( id_4918, id_4913, id_4916);
nand ( id_4976, id_4971, id_4974);
nand ( id_4398, id_4396, id_4397);
nand ( id_4456, id_4454, id_4455);
not ( id_4520, id_4514);
nand ( id_4523, id_4514, id_4521);
not ( id_4608, id_4602);
nand ( id_4611, id_4602, id_4609);
nand ( id_4862, id_4860, id_4861);
nand ( id_4920, id_4918, id_4919);
nand ( id_4978, id_4976, id_4977);
not ( id_5062, id_5056);
nand ( id_5065, id_5056, id_5063);
nand ( id_4522, id_4517, id_4520);
nand ( id_4610, id_4605, id_4608);
nand ( id_5064, id_5059, id_5062);
not ( id_4404, id_4398);
nand ( id_1488, id_4398, id_4405);
not ( id_4462, id_4456);
nand ( id_1493, id_4456, id_4463);
not ( id_4868, id_4862);
nand ( id_2165, id_4862, id_4869);
not ( id_4926, id_4920);
nand ( id_2170, id_4920, id_4927);
nand ( id_4524, id_4522, id_4523);
nand ( id_4612, id_4610, id_4611);
not ( id_4984, id_4978);
nand ( id_4987, id_4978, id_4985);
nand ( id_5066, id_5064, id_5065);
nand ( id_1487, id_4401, id_4404);
nand ( id_1492, id_4459, id_4462);
nand ( id_2164, id_4865, id_4868);
nand ( id_2169, id_4923, id_4926);
nand ( id_4986, id_4981, id_4984);
nand ( id_1489, id_1487, id_1488);
nand ( id_1494, id_1492, id_1493);
nand ( id_2166, id_2164, id_2165);
nand ( id_2171, id_2169, id_2170);
not ( id_4530, id_4524);
nand ( id_4533, id_4524, id_4531);
not ( id_4618, id_4612);
nand ( id_4543, id_4612, id_4619);
nand ( id_4988, id_4986, id_4987);
not ( id_5072, id_5066);
nand ( id_4997, id_5066, id_5073);
nand ( id_4532, id_4527, id_4530);
nand ( id_4542, id_4615, id_4618);
nand ( id_4996, id_5069, id_5072);
and ( id_1513, id_1494, id_1462, id_1502);
and ( id_1514, id_1489, id_1458);
and ( id_1515, id_1494, id_1483);
and ( id_1516, id_1489, id_1486, id_1497);
not ( id_4994, id_4988);
nand ( id_2184, id_4988, id_4995);
and ( id_2190, id_2171, id_2139, id_2179);
and ( id_2191, id_2166, id_2135);
and ( id_2192, id_2171, id_2160);
and ( id_2193, id_2166, id_2163, id_2174);
nand ( id_4534, id_4532, id_4533);
nand ( id_4544, id_4542, id_4543);
nand ( id_4998, id_4996, id_4997);
nand ( id_2183, id_4991, id_4994);
or ( id_4620, id_1513, id_1514, id_1515, id_1516);
or ( id_5074, id_2190, id_2191, id_2192, id_2193);
not ( id_4540, id_4534);
nand ( id_1507, id_4534, id_4541);
not ( id_4550, id_4544);
nand ( id_1510, id_4544, id_4551);
nand ( id_2185, id_2183, id_2184);
not ( id_5004, id_4998);
nand ( id_2187, id_4998, id_5005);
nand ( id_1506, id_4537, id_4540);
nand ( id_1509, id_4547, id_4550);
not ( id_4626, id_4620);
nand ( id_2186, id_5001, id_5004);
and ( id_2195, id_2174, id_2185);
not ( id_5080, id_5074);
nand ( id_1508, id_1506, id_1507);
nand ( id_1511, id_1509, id_1510);
nand ( id_2188, id_2186, id_2187);
not ( id_1512, id_1511);
and ( id_1518, id_1497, id_1508);
not ( id_2189, id_2188);
and ( id_1517, id_1512, id_1502);
and ( id_2194, id_2189, id_2179);
or ( id_4623, id_1517, id_1518);
or ( id_5077, id_2194, id_2195);
nand ( id_1519, id_4623, id_4626);
not ( id_4627, id_4623);
nand ( id_2196, id_5077, id_5080);
not ( id_5081, id_5077);
nand ( id_1520, id_4620, id_4627);
nand ( id_2197, id_5074, id_5081);
nand ( id_1521, id_1519, id_1520);
nand ( id_2198, id_2196, id_2197);
and ( id_840, id_2198, id_3795);
and ( id_879, id_1521, id_3737);
not ( id_1524, id_1521);
not ( id_2201, id_2198);
or ( id_843, id_839, id_840, id_841, id_842);
or ( id_882, id_878, id_879, id_880, id_881);
and ( id_3649, id_1524, id_3628);
and ( id_3652, id_2201, id_3628);
or ( id_3657, id_3648, id_3649);
or ( id_3658, id_3651, id_3652);
and ( id_3636, id_3657, id_3622);
and ( id_3639, id_3658, id_3622);
and ( id_3642, id_3657, id_3622);
and ( id_3645, id_3658, id_3622);
or ( id_3653, id_3636, id_3637);
or ( id_3654, id_3639, id_3640);
or ( id_3655, id_3642, id_3643);
or ( id_3656, id_3645, id_3646);
and ( id_763, id_3656, id_2430, id_2454);
and ( id_764, id_3655, id_2418, id_2454);
and ( id_803, id_3656, id_2488, id_2512);
and ( id_804, id_3655, id_2476, id_2512);
and ( id_1657, id_3654, id_1621, id_1645);
and ( id_1659, id_3653, id_1609, id_1645);
and ( id_2328, id_3654, id_2293, id_2316);
and ( id_2330, id_3653, id_2281, id_2316);
or ( id_1662, id_1657, id_1659, id_1660, id_1661);
or ( id_2333, id_2328, id_2330, id_2331, id_2332);
or ( id_767, id_763, id_764, id_765, id_766);
or ( id_807, id_803, id_804, id_805, id_806);
and ( id_657, id_1662, id_1606);
and ( id_689, id_2333, id_2279);
not ( id_658, id_657);
not ( id_690, id_689);

endmodule
