module c432nr
( id_1gat ,id_4gat ,id_8gat ,id_11gat ,id_14gat ,id_17gat ,id_21gat ,id_24gat ,id_27gat ,id_30gat ,id_34gat ,id_37gat ,id_40gat ,id_43gat ,id_47gat ,id_50gat ,id_53gat ,id_56gat ,id_60gat ,id_63gat ,id_66gat ,id_69gat ,id_73gat ,id_76gat ,id_79gat ,id_82gat ,id_86gat ,id_89gat ,id_92gat ,id_95gat ,id_99gat ,id_102gat ,id_105gat ,id_108gat ,id_112gat ,id_115gat ,id_223gat ,id_329gat ,id_370gat ,id_421gat ,id_430gat ,id_431gat ,id_432gat  );

input id_1gat, id_4gat, id_8gat, id_11gat, id_14gat, id_17gat, id_21gat, id_24gat, id_27gat, id_30gat, id_34gat, id_37gat, id_40gat, id_43gat, id_47gat, id_50gat, id_53gat, id_56gat, id_60gat, id_63gat, id_66gat, id_69gat, id_73gat, id_76gat, id_79gat, id_82gat, id_86gat, id_89gat, id_92gat, id_95gat, id_99gat, id_102gat, id_105gat, id_108gat, id_112gat, id_115gat;

output id_223gat, id_329gat, id_370gat, id_421gat, id_430gat, id_431gat, id_432gat;

not ( id_118gat, id_1gat);
not ( id_119gat, id_4gat);
not ( id_122gat, id_11gat);
not ( id_123gat, id_17gat);
not ( id_126gat, id_24gat);
not ( id_127gat, id_30gat);
not ( id_130gat, id_37gat);
not ( id_131gat, id_43gat);
not ( id_134gat, id_50gat);
not ( id_135gat, id_56gat);
not ( id_138gat, id_63gat);
not ( id_139gat, id_69gat);
not ( id_142gat, id_76gat);
not ( id_143gat, id_82gat);
not ( id_146gat, id_89gat);
not ( id_147gat, id_95gat);
not ( id_150gat, id_102gat);
not ( id_151gat, id_108gat);
nand ( id_154gat, id_118gat, id_4gat);
nor ( id_157gat, id_8gat, id_119gat);
nor ( id_158gat, id_14gat, id_119gat);
nand ( id_159gat, id_122gat, id_17gat);
nand ( id_162gat, id_126gat, id_30gat);
nand ( id_165gat, id_130gat, id_43gat);
nand ( id_168gat, id_134gat, id_56gat);
nand ( id_171gat, id_138gat, id_69gat);
nand ( id_174gat, id_142gat, id_82gat);
nand ( id_177gat, id_146gat, id_95gat);
nand ( id_180gat, id_150gat, id_108gat);
nor ( id_183gat, id_21gat, id_123gat);
nor ( id_184gat, id_27gat, id_123gat);
nor ( id_185gat, id_34gat, id_127gat);
nor ( id_186gat, id_40gat, id_127gat);
nor ( id_187gat, id_47gat, id_131gat);
nor ( id_188gat, id_53gat, id_131gat);
nor ( id_189gat, id_60gat, id_135gat);
nor ( id_190gat, id_66gat, id_135gat);
nor ( id_191gat, id_73gat, id_139gat);
nor ( id_192gat, id_79gat, id_139gat);
nor ( id_193gat, id_86gat, id_143gat);
nor ( id_194gat, id_92gat, id_143gat);
nor ( id_195gat, id_99gat, id_147gat);
nor ( id_196gat, id_105gat, id_147gat);
nor ( id_197gat, id_112gat, id_151gat);
nor ( id_198gat, id_115gat, id_151gat);
and ( id_199gat, id_154gat, id_159gat, id_162gat, id_165gat, id_168gat, id_171gat, id_174gat, id_177gat, id_180gat);
not ( id_203gat, id_199gat);
not ( id_213gat, id_199gat);
not ( id_223gat, id_199gat);
xor ( id_224gat, id_203gat, id_154gat);
xor ( id_227gat, id_203gat, id_159gat);
xor ( id_230gat, id_203gat, id_162gat);
xor ( id_233gat, id_203gat, id_165gat);
xor ( id_236gat, id_203gat, id_168gat);
xor ( id_239gat, id_203gat, id_171gat);
nand ( id_242gat, id_1gat, id_213gat);
xor ( id_243gat, id_203gat, id_174gat);
nand ( id_246gat, id_213gat, id_11gat);
xor ( id_247gat, id_203gat, id_177gat);
nand ( id_250gat, id_213gat, id_24gat);
xor ( id_251gat, id_203gat, id_180gat);
nand ( id_254gat, id_213gat, id_37gat);
nand ( id_255gat, id_213gat, id_50gat);
nand ( id_256gat, id_213gat, id_63gat);
nand ( id_257gat, id_213gat, id_76gat);
nand ( id_258gat, id_213gat, id_89gat);
nand ( id_260gat, id_224gat, id_157gat);
nand ( id_263gat, id_224gat, id_158gat);
nand ( id_264gat, id_227gat, id_183gat);
nand ( id_267gat, id_230gat, id_185gat);
nand ( id_270gat, id_233gat, id_187gat);
nand ( id_273gat, id_236gat, id_189gat);
nand ( id_276gat, id_239gat, id_191gat);
nand ( id_279gat, id_243gat, id_193gat);
nand ( id_282gat, id_247gat, id_195gat);
nand ( id_285gat, id_251gat, id_197gat);
nand ( id_288gat, id_227gat, id_184gat);
nand ( id_289gat, id_230gat, id_186gat);
nand ( id_290gat, id_233gat, id_188gat);
nand ( id_291gat, id_236gat, id_190gat);
nand ( id_292gat, id_239gat, id_192gat);
nand ( id_293gat, id_243gat, id_194gat);
nand ( id_294gat, id_247gat, id_196gat);
nand ( id_295gat, id_251gat, id_198gat);
and ( id_296gat, id_260gat, id_264gat, id_267gat, id_270gat, id_273gat, id_276gat, id_279gat, id_282gat, id_285gat);
not ( id_300gat, id_263gat);
not ( id_301gat, id_288gat);
not ( id_302gat, id_289gat);
not ( id_303gat, id_290gat);
not ( id_304gat, id_291gat);
not ( id_305gat, id_292gat);
not ( id_306gat, id_293gat);
not ( id_307gat, id_294gat);
not ( id_308gat, id_295gat);
not ( id_309gat, id_296gat);
not ( id_319gat, id_296gat);
not ( id_329gat, id_296gat);
xor ( id_330gat, id_309gat, id_260gat);
xor ( id_331gat, id_309gat, id_264gat);
xor ( id_332gat, id_309gat, id_267gat);
xor ( id_333gat, id_309gat, id_270gat);
nand ( id_334gat, id_8gat, id_319gat);
xor ( id_335gat, id_309gat, id_273gat);
nand ( id_336gat, id_319gat, id_21gat);
xor ( id_337gat, id_309gat, id_276gat);
nand ( id_338gat, id_319gat, id_34gat);
xor ( id_339gat, id_309gat, id_279gat);
nand ( id_340gat, id_319gat, id_47gat);
xor ( id_341gat, id_309gat, id_282gat);
nand ( id_342gat, id_319gat, id_60gat);
xor ( id_343gat, id_309gat, id_285gat);
nand ( id_344gat, id_319gat, id_73gat);
nand ( id_345gat, id_319gat, id_86gat);
nand ( id_346gat, id_319gat, id_99gat);
nand ( id_348gat, id_330gat, id_300gat);
nand ( id_349gat, id_331gat, id_301gat);
nand ( id_350gat, id_332gat, id_302gat);
nand ( id_351gat, id_333gat, id_303gat);
nand ( id_352gat, id_335gat, id_304gat);
nand ( id_353gat, id_337gat, id_305gat);
nand ( id_354gat, id_339gat, id_306gat);
nand ( id_355gat, id_341gat, id_307gat);
nand ( id_356gat, id_343gat, id_308gat);
and ( id_357gat, id_348gat, id_349gat, id_350gat, id_351gat, id_352gat, id_353gat, id_354gat, id_355gat, id_356gat);
not ( id_360gat, id_357gat);
not ( id_370gat, id_357gat);
nand ( id_371gat, id_14gat, id_360gat);
nand ( id_372gat, id_360gat, id_27gat);
nand ( id_373gat, id_360gat, id_40gat);
nand ( id_374gat, id_360gat, id_53gat);
nand ( id_375gat, id_360gat, id_66gat);
nand ( id_376gat, id_360gat, id_79gat);
nand ( id_377gat, id_360gat, id_92gat);
nand ( id_378gat, id_360gat, id_105gat);
nand ( id_380gat, id_4gat, id_242gat, id_334gat, id_371gat);
nand ( id_381gat, id_246gat, id_336gat, id_372gat, id_17gat);
nand ( id_386gat, id_250gat, id_338gat, id_373gat, id_30gat);
nand ( id_393gat, id_254gat, id_340gat, id_374gat, id_43gat);
nand ( id_399gat, id_255gat, id_342gat, id_375gat, id_56gat);
nand ( id_404gat, id_256gat, id_344gat, id_376gat, id_69gat);
nand ( id_407gat, id_257gat, id_345gat, id_377gat, id_82gat);
nand ( id_411gat, id_258gat, id_346gat, id_378gat, id_95gat);
not ( id_414gat, id_108gat);
not ( id_415gat, id_380gat);
and ( id_416gat, id_381gat, id_386gat, id_393gat, id_399gat, id_404gat, id_407gat, id_411gat, id_414gat);
not ( id_417gat, id_393gat);
not ( id_418gat, id_404gat);
not ( id_419gat, id_407gat);
not ( id_420gat, id_411gat);
nor ( id_421gat, id_415gat, id_416gat);
nand ( id_422gat, id_386gat, id_417gat);
nand ( id_425gat, id_386gat, id_393gat, id_418gat, id_399gat);
nand ( id_428gat, id_399gat, id_393gat, id_419gat);
nand ( id_429gat, id_386gat, id_407gat, id_420gat);
nand ( id_430gat, id_381gat, id_386gat, id_422gat, id_399gat);
nand ( id_431gat, id_381gat, id_386gat, id_425gat, id_428gat);
nand ( id_432gat, id_381gat, id_422gat, id_425gat, id_429gat);

endmodule
