module c499nr
( id_id0 ,id_id1 ,id_id2 ,id_id3 ,id_id4 ,id_id5 ,id_id6 ,id_id7 ,id_id8 ,id_id9 ,id_id10 ,id_id11 ,id_id12 ,id_id13 ,id_id14 ,id_id15 ,id_id16 ,id_id17 ,id_id18 ,id_id19 ,id_id20 ,id_id21 ,id_id22 ,id_id23 ,id_id24 ,id_id25 ,id_id26 ,id_id27 ,id_id28 ,id_id29 ,id_id30 ,id_id31 ,id_ic0 ,id_ic1 ,id_ic2 ,id_ic3 ,id_ic4 ,id_ic5 ,id_ic6 ,id_ic7 ,id_r ,id_od0 ,id_od1 ,id_od2 ,id_od3 ,id_od4 ,id_od5 ,id_od6 ,id_od7 ,id_od8 ,id_od9 ,id_od10 ,id_od11 ,id_od12 ,id_od13 ,id_od14 ,id_od15 ,id_od16 ,id_od17 ,id_od18 ,id_od19 ,id_od20 ,id_od21 ,id_od22 ,id_od23 ,id_od24 ,id_od25 ,id_od26 ,id_od27 ,id_od28 ,id_od29 ,id_od30 ,id_od31  );

input id_id0, id_id1, id_id2, id_id3, id_id4, id_id5, id_id6, id_id7, id_id8, id_id9, id_id10, id_id11, id_id12, id_id13, id_id14, id_id15, id_id16, id_id17, id_id18, id_id19, id_id20, id_id21, id_id22, id_id23, id_id24, id_id25, id_id26, id_id27, id_id28, id_id29, id_id30, id_id31, id_ic0, id_ic1, id_ic2, id_ic3, id_ic4, id_ic5, id_ic6, id_ic7, id_r;

output id_od0, id_od1, id_od2, id_od3, id_od4, id_od5, id_od6, id_od7, id_od8, id_od9, id_od10, id_od11, id_od12, id_od13, id_od14, id_od15, id_od16, id_od17, id_od18, id_od19, id_od20, id_od21, id_od22, id_od23, id_od24, id_od25, id_od26, id_od27, id_od28, id_od29, id_od30, id_od31;

xor ( id_xa0, id_id0, id_id1);
xor ( id_xa1, id_id2, id_id3);
xor ( id_xa2, id_id4, id_id5);
xor ( id_xa3, id_id6, id_id7);
xor ( id_xa4, id_id8, id_id9);
xor ( id_xa5, id_id10, id_id11);
xor ( id_xa6, id_id12, id_id13);
xor ( id_xa7, id_id14, id_id15);
xor ( id_xa8, id_id16, id_id17);
xor ( id_xa9, id_id18, id_id19);
xor ( id_xa10, id_id20, id_id21);
xor ( id_xa11, id_id22, id_id23);
xor ( id_xa12, id_id24, id_id25);
xor ( id_xa13, id_id26, id_id27);
xor ( id_xa14, id_id28, id_id29);
xor ( id_xa15, id_id30, id_id31);
and ( id_h0, id_ic0, id_r);
and ( id_h1, id_ic1, id_r);
and ( id_h2, id_ic2, id_r);
and ( id_h3, id_ic3, id_r);
and ( id_h4, id_ic4, id_r);
and ( id_h5, id_ic5, id_r);
and ( id_h6, id_ic6, id_r);
and ( id_h7, id_ic7, id_r);
xor ( id_xb0, id_id0, id_id4);
xor ( id_xc0, id_id8, id_id12);
xor ( id_xb1, id_id1, id_id5);
xor ( id_xc1, id_id9, id_id13);
xor ( id_xb2, id_id2, id_id6);
xor ( id_xc2, id_id10, id_id14);
xor ( id_xb3, id_id3, id_id7);
xor ( id_xc3, id_id11, id_id15);
xor ( id_xb4, id_id16, id_id20);
xor ( id_xc4, id_id24, id_id28);
xor ( id_xb5, id_id17, id_id21);
xor ( id_xc5, id_id25, id_id29);
xor ( id_xb6, id_id18, id_id22);
xor ( id_xc6, id_id26, id_id30);
xor ( id_xb7, id_id19, id_id23);
xor ( id_xc7, id_id27, id_id31);
xor ( id_f0, id_xa0, id_xa1);
xor ( id_f1, id_xa2, id_xa3);
xor ( id_f2, id_xa4, id_xa5);
xor ( id_f3, id_xa6, id_xa7);
xor ( id_f4, id_xa8, id_xa9);
xor ( id_f5, id_xa10, id_xa11);
xor ( id_f6, id_xa12, id_xa13);
xor ( id_f7, id_xa14, id_xa15);
xor ( id_xe0, id_xb0, id_xc0);
xor ( id_xe1, id_xb1, id_xc1);
xor ( id_xe2, id_xb2, id_xc2);
xor ( id_xe3, id_xb3, id_xc3);
xor ( id_xe4, id_xb4, id_xc4);
xor ( id_xe5, id_xb5, id_xc5);
xor ( id_xe6, id_xb6, id_xc6);
xor ( id_xe7, id_xb7, id_xc7);
xor ( id_g0, id_f0, id_f1);
xor ( id_g1, id_f2, id_f3);
xor ( id_g2, id_f0, id_f2);
xor ( id_g3, id_f1, id_f3);
xor ( id_g4, id_f4, id_f5);
xor ( id_g5, id_f6, id_f7);
xor ( id_g6, id_f4, id_f6);
xor ( id_g7, id_f5, id_f7);
xor ( id_xd0, id_h0, id_g4);
xor ( id_xd1, id_h1, id_g5);
xor ( id_xd2, id_h2, id_g6);
xor ( id_xd3, id_h3, id_g7);
xor ( id_xd4, id_h4, id_g0);
xor ( id_xd5, id_h5, id_g1);
xor ( id_xd6, id_h6, id_g2);
xor ( id_xd7, id_h7, id_g3);
xor ( id_s0, id_xe0, id_xd0);
xor ( id_s1, id_xe1, id_xd1);
xor ( id_s2, id_xe2, id_xd2);
xor ( id_s3, id_xe3, id_xd3);
xor ( id_s4, id_xe4, id_xd4);
xor ( id_s5, id_xe5, id_xd5);
xor ( id_s6, id_xe6, id_xd6);
xor ( id_s7, id_xe7, id_xd7);
not ( id_y0a, id_s0);
not ( id_y1a, id_s1);
not ( id_y2a, id_s2);
not ( id_y0b, id_s0);
not ( id_y1b, id_s1);
not ( id_y3b, id_s3);
not ( id_y0c, id_s0);
not ( id_y2c, id_s2);
not ( id_y3c, id_s3);
not ( id_y1d, id_s1);
not ( id_y2d, id_s2);
not ( id_y3d, id_s3);
not ( id_y5i, id_s5);
not ( id_y7i, id_s7);
not ( id_y5j, id_s5);
not ( id_y6j, id_s6);
not ( id_y4k, id_s4);
not ( id_y7k, id_s7);
not ( id_y4l, id_s4);
not ( id_y6l, id_s6);
not ( id_y4a, id_s4);
not ( id_y5a, id_s5);
not ( id_y6a, id_s6);
not ( id_y4b, id_s4);
not ( id_y5b, id_s5);
not ( id_y7b, id_s7);
not ( id_y4c, id_s4);
not ( id_y6c, id_s6);
not ( id_y7c, id_s7);
not ( id_y5d, id_s5);
not ( id_y6d, id_s6);
not ( id_y7d, id_s7);
not ( id_y1i, id_s1);
not ( id_y3i, id_s3);
not ( id_y1j, id_s1);
not ( id_y2j, id_s2);
not ( id_y0k, id_s0);
not ( id_y3k, id_s3);
not ( id_y0l, id_s0);
not ( id_y2l, id_s2);
and ( id_t0, id_y0a, id_y1a, id_y2a);
and ( id_t1, id_y0b, id_y1b, id_y3b);
and ( id_t2, id_y0c, id_y2c, id_y3c);
and ( id_t3, id_y1d, id_y2d, id_y3d);
and ( id_t4, id_y4a, id_y5a, id_y6a);
and ( id_t5, id_y4b, id_y5b, id_y7b);
and ( id_t6, id_y4c, id_y6c, id_y7c);
and ( id_t7, id_y5d, id_y6d, id_y7d);
or ( id_u0, id_t0, id_t1, id_t2, id_t3);
or ( id_u1, id_t4, id_t5, id_t6, id_t7);
and ( id_wa, id_s4, id_y5i, id_s6, id_y7i, id_u0);
and ( id_wb, id_s4, id_y5j, id_y6j, id_s7, id_u0);
and ( id_wc, id_y4k, id_s5, id_s6, id_y7k, id_u0);
and ( id_wd, id_y4l, id_s5, id_y6l, id_s7, id_u0);
and ( id_we, id_s0, id_y1i, id_s2, id_y3i, id_u1);
and ( id_wf, id_s0, id_y1j, id_y2j, id_s3, id_u1);
and ( id_wg, id_y0k, id_s1, id_s2, id_y3k, id_u1);
and ( id_wh, id_y0l, id_s1, id_y2l, id_s3, id_u1);
and ( id_e0, id_s0, id_wa);
and ( id_e1, id_s1, id_wa);
and ( id_e2, id_s2, id_wa);
and ( id_e3, id_s3, id_wa);
and ( id_e4, id_s0, id_wb);
and ( id_e5, id_s1, id_wb);
and ( id_e6, id_s2, id_wb);
and ( id_e7, id_s3, id_wb);
and ( id_e8, id_s0, id_wc);
and ( id_e9, id_s1, id_wc);
and ( id_e10, id_s2, id_wc);
and ( id_e11, id_s3, id_wc);
and ( id_e12, id_s0, id_wd);
and ( id_e13, id_s1, id_wd);
and ( id_e14, id_s2, id_wd);
and ( id_e15, id_s3, id_wd);
and ( id_e16, id_s4, id_we);
and ( id_e17, id_s5, id_we);
and ( id_e18, id_s6, id_we);
and ( id_e19, id_s7, id_we);
and ( id_e20, id_s4, id_wf);
and ( id_e21, id_s5, id_wf);
and ( id_e22, id_s6, id_wf);
and ( id_e23, id_s7, id_wf);
and ( id_e24, id_s4, id_wg);
and ( id_e25, id_s5, id_wg);
and ( id_e26, id_s6, id_wg);
and ( id_e27, id_s7, id_wg);
and ( id_e28, id_s4, id_wh);
and ( id_e29, id_s5, id_wh);
and ( id_e30, id_s6, id_wh);
and ( id_e31, id_s7, id_wh);
xor ( id_od0, id_id0, id_e0);
xor ( id_od1, id_id1, id_e1);
xor ( id_od2, id_id2, id_e2);
xor ( id_od3, id_id3, id_e3);
xor ( id_od4, id_id4, id_e4);
xor ( id_od5, id_id5, id_e5);
xor ( id_od6, id_id6, id_e6);
xor ( id_od7, id_id7, id_e7);
xor ( id_od8, id_id8, id_e8);
xor ( id_od9, id_id9, id_e9);
xor ( id_od10, id_id10, id_e10);
xor ( id_od11, id_id11, id_e11);
xor ( id_od12, id_id12, id_e12);
xor ( id_od13, id_id13, id_e13);
xor ( id_od14, id_id14, id_e14);
xor ( id_od15, id_id15, id_e15);
xor ( id_od16, id_id16, id_e16);
xor ( id_od17, id_id17, id_e17);
xor ( id_od18, id_id18, id_e18);
xor ( id_od19, id_id19, id_e19);
xor ( id_od20, id_id20, id_e20);
xor ( id_od21, id_id21, id_e21);
xor ( id_od22, id_id22, id_e22);
xor ( id_od23, id_id23, id_e23);
xor ( id_od24, id_id24, id_e24);
xor ( id_od25, id_id25, id_e25);
xor ( id_od26, id_id26, id_e26);
xor ( id_od27, id_id27, id_e27);
xor ( id_od28, id_id28, id_e28);
xor ( id_od29, id_id29, id_e29);
xor ( id_od30, id_id30, id_e30);
xor ( id_od31, id_id31, id_e31);

endmodule
