module c880
( id_1gat ,id_8gat ,id_13gat ,id_17gat ,id_26gat ,id_29gat ,id_36gat ,id_42gat ,id_51gat ,id_55gat ,id_59gat ,id_68gat ,id_72gat ,id_73gat ,id_74gat ,id_75gat ,id_80gat ,id_85gat ,id_86gat ,id_87gat ,id_88gat ,id_89gat ,id_90gat ,id_91gat ,id_96gat ,id_101gat ,id_106gat ,id_111gat ,id_116gat ,id_121gat ,id_126gat ,id_130gat ,id_135gat ,id_138gat ,id_143gat ,id_146gat ,id_149gat ,id_152gat ,id_153gat ,id_156gat ,id_159gat ,id_165gat ,id_171gat ,id_177gat ,id_183gat ,id_189gat ,id_195gat ,id_201gat ,id_207gat ,id_210gat ,id_219gat ,id_228gat ,id_237gat ,id_246gat ,id_255gat ,id_259gat ,id_260gat ,id_261gat ,id_267gat ,id_268gat ,id_388gat ,id_389gat ,id_390gat ,id_391gat ,id_418gat ,id_419gat ,id_420gat ,id_421gat ,id_422gat ,id_423gat ,id_446gat ,id_447gat ,id_448gat ,id_449gat ,id_450gat ,id_767gat ,id_768gat ,id_850gat ,id_863gat ,id_864gat ,id_865gat ,id_866gat ,id_874gat ,id_878gat ,id_879gat ,id_880gat );

input id_1gat, id_8gat, id_13gat, id_17gat, id_26gat, id_29gat, id_36gat, id_42gat, id_51gat, id_55gat, id_59gat, id_68gat, id_72gat, id_73gat, id_74gat, id_75gat, id_80gat, id_85gat, id_86gat, id_87gat, id_88gat, id_89gat, id_90gat, id_91gat, id_96gat, id_101gat, id_106gat, id_111gat, id_116gat, id_121gat, id_126gat, id_130gat, id_135gat, id_138gat, id_143gat, id_146gat, id_149gat, id_152gat, id_153gat, id_156gat, id_159gat, id_165gat, id_171gat, id_177gat, id_183gat, id_189gat, id_195gat, id_201gat, id_207gat, id_210gat, id_219gat, id_228gat, id_237gat, id_246gat, id_255gat, id_259gat, id_260gat, id_261gat, id_267gat, id_268gat;

output id_388gat, id_389gat, id_390gat, id_391gat, id_418gat, id_419gat, id_420gat, id_421gat, id_422gat, id_423gat, id_446gat, id_447gat, id_448gat, id_449gat, id_450gat, id_767gat, id_768gat, id_850gat, id_863gat, id_864gat, id_865gat, id_866gat, id_874gat, id_878gat, id_879gat, id_880gat;

nand ( id_269gat, id_1gat, id_8gat, id_13gat, id_17gat);
nand ( id_270gat, id_1gat, id_26gat, id_13gat, id_17gat);
and ( id_273gat, id_29gat, id_36gat, id_42gat);
and ( id_276gat, id_1gat, id_26gat, id_51gat);
nand ( id_279gat, id_1gat, id_8gat, id_51gat, id_17gat);
nand ( id_280gat, id_1gat, id_8gat, id_13gat, id_55gat);
nand ( id_284gat, id_59gat, id_42gat, id_68gat, id_72gat);
nand ( id_285gat, id_29gat, id_68gat);
nand ( id_286gat, id_59gat, id_68gat, id_74gat);
and ( id_287gat, id_29gat, id_75gat, id_80gat);
and ( id_290gat, id_29gat, id_75gat, id_42gat);
and ( id_291gat, id_29gat, id_36gat, id_80gat);
and ( id_292gat, id_29gat, id_36gat, id_42gat);
and ( id_293gat, id_59gat, id_75gat, id_80gat);
and ( id_294gat, id_59gat, id_75gat, id_42gat);
and ( id_295gat, id_59gat, id_36gat, id_80gat);
and ( id_296gat, id_59gat, id_36gat, id_42gat);
and ( id_297gat, id_85gat, id_86gat);
or ( id_298gat, id_87gat, id_88gat);
nand ( id_301gat, id_91gat, id_96gat);
or ( id_302gat, id_91gat, id_96gat);
nand ( id_303gat, id_101gat, id_106gat);
or ( id_304gat, id_101gat, id_106gat);
nand ( id_305gat, id_111gat, id_116gat);
or ( id_306gat, id_111gat, id_116gat);
nand ( id_307gat, id_121gat, id_126gat);
or ( id_308gat, id_121gat, id_126gat);
and ( id_309gat, id_8gat, id_138gat);
not ( id_310gat, id_268gat);
and ( id_316gat, id_51gat, id_138gat);
and ( id_317gat, id_17gat, id_138gat);
and ( id_318gat, id_152gat, id_138gat);
nand ( id_319gat, id_59gat, id_156gat);
nor ( id_322gat, id_17gat, id_42gat);
and ( id_323gat, id_17gat, id_42gat);
nand ( id_324gat, id_159gat, id_165gat);
or ( id_325gat, id_159gat, id_165gat);
nand ( id_326gat, id_171gat, id_177gat);
or ( id_327gat, id_171gat, id_177gat);
nand ( id_328gat, id_183gat, id_189gat);
or ( id_329gat, id_183gat, id_189gat);
nand ( id_330gat, id_195gat, id_201gat);
or ( id_331gat, id_195gat, id_201gat);
and ( id_332gat, id_210gat, id_91gat);
and ( id_333gat, id_210gat, id_96gat);
and ( id_334gat, id_210gat, id_101gat);
and ( id_335gat, id_210gat, id_106gat);
and ( id_336gat, id_210gat, id_111gat);
and ( id_337gat, id_255gat, id_259gat);
and ( id_338gat, id_210gat, id_116gat);
and ( id_339gat, id_255gat, id_260gat);
and ( id_340gat, id_210gat, id_121gat);
and ( id_341gat, id_255gat, id_267gat);
not ( id_342gat, id_269gat);
not ( id_343gat, id_273gat);
or ( id_344gat, id_270gat, id_273gat);
not ( id_345gat, id_276gat);
not ( id_346gat, id_276gat);
not ( id_347gat, id_279gat);
nor ( id_348gat, id_280gat, id_284gat);
or ( id_349gat, id_280gat, id_285gat);
or ( id_350gat, id_280gat, id_286gat);
not ( id_351gat, id_293gat);
not ( id_352gat, id_294gat);
not ( id_353gat, id_295gat);
not ( id_354gat, id_296gat);
nand ( id_355gat, id_89gat, id_298gat);
and ( id_356gat, id_90gat, id_298gat);
nand ( id_357gat, id_301gat, id_302gat);
nand ( id_360gat, id_303gat, id_304gat);
nand ( id_363gat, id_305gat, id_306gat);
nand ( id_366gat, id_307gat, id_308gat);
not ( id_369gat, id_310gat);
nor ( id_375gat, id_322gat, id_323gat);
nand ( id_376gat, id_324gat, id_325gat);
nand ( id_379gat, id_326gat, id_327gat);
nand ( id_382gat, id_328gat, id_329gat);
nand ( id_385gat, id_330gat, id_331gat);
buf ( id_388gat, id_290gat);
buf ( id_389gat, id_291gat);
buf ( id_390gat, id_292gat);
buf ( id_391gat, id_297gat);
or ( id_392gat, id_270gat, id_343gat);
not ( id_393gat, id_345gat);
not ( id_399gat, id_346gat);
and ( id_400gat, id_348gat, id_73gat);
not ( id_401gat, id_349gat);
not ( id_402gat, id_350gat);
not ( id_403gat, id_355gat);
not ( id_404gat, id_357gat);
not ( id_405gat, id_360gat);
and ( id_406gat, id_357gat, id_360gat);
not ( id_407gat, id_363gat);
not ( id_408gat, id_366gat);
and ( id_409gat, id_363gat, id_366gat);
nand ( id_410gat, id_347gat, id_352gat);
not ( id_411gat, id_376gat);
not ( id_412gat, id_379gat);
and ( id_413gat, id_376gat, id_379gat);
not ( id_414gat, id_382gat);
not ( id_415gat, id_385gat);
and ( id_416gat, id_382gat, id_385gat);
and ( id_417gat, id_210gat, id_369gat);
buf ( id_418gat, id_342gat);
buf ( id_419gat, id_344gat);
buf ( id_420gat, id_351gat);
buf ( id_421gat, id_353gat);
buf ( id_422gat, id_354gat);
buf ( id_423gat, id_356gat);
not ( id_424gat, id_400gat);
and ( id_425gat, id_404gat, id_405gat);
and ( id_426gat, id_407gat, id_408gat);
and ( id_427gat, id_319gat, id_393gat, id_55gat);
and ( id_432gat, id_393gat, id_17gat, id_287gat);
nand ( id_437gat, id_393gat, id_287gat, id_55gat);
nand ( id_442gat, id_375gat, id_59gat, id_156gat, id_393gat);
nand ( id_443gat, id_393gat, id_319gat, id_17gat);
and ( id_444gat, id_411gat, id_412gat);
and ( id_445gat, id_414gat, id_415gat);
buf ( id_446gat, id_392gat);
buf ( id_447gat, id_399gat);
buf ( id_448gat, id_401gat);
buf ( id_449gat, id_402gat);
buf ( id_450gat, id_403gat);
not ( id_451gat, id_424gat);
nor ( id_460gat, id_406gat, id_425gat);
nor ( id_463gat, id_409gat, id_426gat);
nand ( id_466gat, id_442gat, id_410gat);
and ( id_475gat, id_143gat, id_427gat);
and ( id_476gat, id_310gat, id_432gat);
and ( id_477gat, id_146gat, id_427gat);
and ( id_478gat, id_310gat, id_432gat);
and ( id_479gat, id_149gat, id_427gat);
and ( id_480gat, id_310gat, id_432gat);
and ( id_481gat, id_153gat, id_427gat);
and ( id_482gat, id_310gat, id_432gat);
nand ( id_483gat, id_443gat, id_1gat);
or ( id_488gat, id_369gat, id_437gat);
or ( id_489gat, id_369gat, id_437gat);
or ( id_490gat, id_369gat, id_437gat);
or ( id_491gat, id_369gat, id_437gat);
nor ( id_492gat, id_413gat, id_444gat);
nor ( id_495gat, id_416gat, id_445gat);
nand ( id_498gat, id_130gat, id_460gat);
or ( id_499gat, id_130gat, id_460gat);
nand ( id_500gat, id_463gat, id_135gat);
or ( id_501gat, id_463gat, id_135gat);
and ( id_502gat, id_91gat, id_466gat);
nor ( id_503gat, id_475gat, id_476gat);
and ( id_504gat, id_96gat, id_466gat);
nor ( id_505gat, id_477gat, id_478gat);
and ( id_506gat, id_101gat, id_466gat);
nor ( id_507gat, id_479gat, id_480gat);
and ( id_508gat, id_106gat, id_466gat);
nor ( id_509gat, id_481gat, id_482gat);
and ( id_510gat, id_143gat, id_483gat);
and ( id_511gat, id_111gat, id_466gat);
and ( id_512gat, id_146gat, id_483gat);
and ( id_513gat, id_116gat, id_466gat);
and ( id_514gat, id_149gat, id_483gat);
and ( id_515gat, id_121gat, id_466gat);
and ( id_516gat, id_153gat, id_483gat);
and ( id_517gat, id_126gat, id_466gat);
nand ( id_518gat, id_130gat, id_492gat);
or ( id_519gat, id_130gat, id_492gat);
nand ( id_520gat, id_495gat, id_207gat);
or ( id_521gat, id_495gat, id_207gat);
and ( id_522gat, id_451gat, id_159gat);
and ( id_523gat, id_451gat, id_165gat);
and ( id_524gat, id_451gat, id_171gat);
and ( id_525gat, id_451gat, id_177gat);
and ( id_526gat, id_451gat, id_183gat);
nand ( id_527gat, id_451gat, id_189gat);
nand ( id_528gat, id_451gat, id_195gat);
nand ( id_529gat, id_451gat, id_201gat);
nand ( id_530gat, id_498gat, id_499gat);
nand ( id_533gat, id_500gat, id_501gat);
nor ( id_536gat, id_309gat, id_502gat);
nor ( id_537gat, id_316gat, id_504gat);
nor ( id_538gat, id_317gat, id_506gat);
nor ( id_539gat, id_318gat, id_508gat);
nor ( id_540gat, id_510gat, id_511gat);
nor ( id_541gat, id_512gat, id_513gat);
nor ( id_542gat, id_514gat, id_515gat);
nor ( id_543gat, id_516gat, id_517gat);
nand ( id_544gat, id_518gat, id_519gat);
nand ( id_547gat, id_520gat, id_521gat);
not ( id_550gat, id_530gat);
not ( id_551gat, id_533gat);
and ( id_552gat, id_530gat, id_533gat);
nand ( id_553gat, id_536gat, id_503gat);
nand ( id_557gat, id_537gat, id_505gat);
nand ( id_561gat, id_538gat, id_507gat);
nand ( id_565gat, id_539gat, id_509gat);
nand ( id_569gat, id_488gat, id_540gat);
nand ( id_573gat, id_489gat, id_541gat);
nand ( id_577gat, id_490gat, id_542gat);
nand ( id_581gat, id_491gat, id_543gat);
not ( id_585gat, id_544gat);
not ( id_586gat, id_547gat);
and ( id_587gat, id_544gat, id_547gat);
and ( id_588gat, id_550gat, id_551gat);
and ( id_589gat, id_585gat, id_586gat);
nand ( id_590gat, id_553gat, id_159gat);
or ( id_593gat, id_553gat, id_159gat);
and ( id_596gat, id_246gat, id_553gat);
nand ( id_597gat, id_557gat, id_165gat);
or ( id_600gat, id_557gat, id_165gat);
and ( id_605gat, id_246gat, id_557gat);
nand ( id_606gat, id_561gat, id_171gat);
or ( id_609gat, id_561gat, id_171gat);
and ( id_615gat, id_246gat, id_561gat);
nand ( id_616gat, id_565gat, id_177gat);
or ( id_619gat, id_565gat, id_177gat);
and ( id_624gat, id_246gat, id_565gat);
nand ( id_625gat, id_569gat, id_183gat);
or ( id_628gat, id_569gat, id_183gat);
and ( id_631gat, id_246gat, id_569gat);
nand ( id_632gat, id_573gat, id_189gat);
or ( id_635gat, id_573gat, id_189gat);
and ( id_640gat, id_246gat, id_573gat);
nand ( id_641gat, id_577gat, id_195gat);
or ( id_644gat, id_577gat, id_195gat);
and ( id_650gat, id_246gat, id_577gat);
nand ( id_651gat, id_581gat, id_201gat);
or ( id_654gat, id_581gat, id_201gat);
and ( id_659gat, id_246gat, id_581gat);
nor ( id_660gat, id_552gat, id_588gat);
nor ( id_661gat, id_587gat, id_589gat);
not ( id_662gat, id_590gat);
and ( id_665gat, id_593gat, id_590gat);
nor ( id_669gat, id_596gat, id_522gat);
not ( id_670gat, id_597gat);
and ( id_673gat, id_600gat, id_597gat);
nor ( id_677gat, id_605gat, id_523gat);
not ( id_678gat, id_606gat);
and ( id_682gat, id_609gat, id_606gat);
nor ( id_686gat, id_615gat, id_524gat);
not ( id_687gat, id_616gat);
and ( id_692gat, id_619gat, id_616gat);
nor ( id_696gat, id_624gat, id_525gat);
not ( id_697gat, id_625gat);
and ( id_700gat, id_628gat, id_625gat);
nor ( id_704gat, id_631gat, id_526gat);
not ( id_705gat, id_632gat);
and ( id_708gat, id_635gat, id_632gat);
nor ( id_712gat, id_337gat, id_640gat);
not ( id_713gat, id_641gat);
and ( id_717gat, id_644gat, id_641gat);
nor ( id_721gat, id_339gat, id_650gat);
not ( id_722gat, id_651gat);
and ( id_727gat, id_654gat, id_651gat);
nor ( id_731gat, id_341gat, id_659gat);
nand ( id_732gat, id_654gat, id_261gat);
nand ( id_733gat, id_644gat, id_654gat, id_261gat);
nand ( id_734gat, id_635gat, id_644gat, id_654gat, id_261gat);
not ( id_735gat, id_662gat);
and ( id_736gat, id_228gat, id_665gat);
and ( id_737gat, id_237gat, id_662gat);
not ( id_738gat, id_670gat);
and ( id_739gat, id_228gat, id_673gat);
and ( id_740gat, id_237gat, id_670gat);
not ( id_741gat, id_678gat);
and ( id_742gat, id_228gat, id_682gat);
and ( id_743gat, id_237gat, id_678gat);
not ( id_744gat, id_687gat);
and ( id_745gat, id_228gat, id_692gat);
and ( id_746gat, id_237gat, id_687gat);
not ( id_747gat, id_697gat);
and ( id_748gat, id_228gat, id_700gat);
and ( id_749gat, id_237gat, id_697gat);
not ( id_750gat, id_705gat);
and ( id_751gat, id_228gat, id_708gat);
and ( id_752gat, id_237gat, id_705gat);
not ( id_753gat, id_713gat);
and ( id_754gat, id_228gat, id_717gat);
and ( id_755gat, id_237gat, id_713gat);
not ( id_756gat, id_722gat);
nor ( id_757gat, id_727gat, id_261gat);
and ( id_758gat, id_727gat, id_261gat);
and ( id_759gat, id_228gat, id_727gat);
and ( id_760gat, id_237gat, id_722gat);
nand ( id_761gat, id_644gat, id_722gat);
nand ( id_762gat, id_635gat, id_713gat);
nand ( id_763gat, id_635gat, id_644gat, id_722gat);
nand ( id_764gat, id_609gat, id_687gat);
nand ( id_765gat, id_600gat, id_678gat);
nand ( id_766gat, id_600gat, id_609gat, id_687gat);
buf ( id_767gat, id_660gat);
buf ( id_768gat, id_661gat);
nor ( id_769gat, id_736gat, id_737gat);
nor ( id_770gat, id_739gat, id_740gat);
nor ( id_771gat, id_742gat, id_743gat);
nor ( id_772gat, id_745gat, id_746gat);
nand ( id_773gat, id_750gat, id_762gat, id_763gat, id_734gat);
nor ( id_777gat, id_748gat, id_749gat);
nand ( id_778gat, id_753gat, id_761gat, id_733gat);
nor ( id_781gat, id_751gat, id_752gat);
nand ( id_782gat, id_756gat, id_732gat);
nor ( id_785gat, id_754gat, id_755gat);
nor ( id_786gat, id_757gat, id_758gat);
nor ( id_787gat, id_759gat, id_760gat);
nor ( id_788gat, id_700gat, id_773gat);
and ( id_789gat, id_700gat, id_773gat);
nor ( id_790gat, id_708gat, id_778gat);
and ( id_791gat, id_708gat, id_778gat);
nor ( id_792gat, id_717gat, id_782gat);
and ( id_793gat, id_717gat, id_782gat);
and ( id_794gat, id_219gat, id_786gat);
nand ( id_795gat, id_628gat, id_773gat);
nand ( id_796gat, id_795gat, id_747gat);
nor ( id_802gat, id_788gat, id_789gat);
nor ( id_803gat, id_790gat, id_791gat);
nor ( id_804gat, id_792gat, id_793gat);
nor ( id_805gat, id_340gat, id_794gat);
nor ( id_806gat, id_692gat, id_796gat);
and ( id_807gat, id_692gat, id_796gat);
and ( id_808gat, id_219gat, id_802gat);
and ( id_809gat, id_219gat, id_803gat);
and ( id_810gat, id_219gat, id_804gat);
nand ( id_811gat, id_805gat, id_787gat, id_731gat, id_529gat);
nand ( id_812gat, id_619gat, id_796gat);
nand ( id_813gat, id_609gat, id_619gat, id_796gat);
nand ( id_814gat, id_600gat, id_609gat, id_619gat, id_796gat);
nand ( id_815gat, id_738gat, id_765gat, id_766gat, id_814gat);
nand ( id_819gat, id_741gat, id_764gat, id_813gat);
nand ( id_822gat, id_744gat, id_812gat);
nor ( id_825gat, id_806gat, id_807gat);
nor ( id_826gat, id_335gat, id_808gat);
nor ( id_827gat, id_336gat, id_809gat);
nor ( id_828gat, id_338gat, id_810gat);
not ( id_829gat, id_811gat);
nor ( id_830gat, id_665gat, id_815gat);
and ( id_831gat, id_665gat, id_815gat);
nor ( id_832gat, id_673gat, id_819gat);
and ( id_833gat, id_673gat, id_819gat);
nor ( id_834gat, id_682gat, id_822gat);
and ( id_835gat, id_682gat, id_822gat);
and ( id_836gat, id_219gat, id_825gat);
nand ( id_837gat, id_826gat, id_777gat, id_704gat);
nand ( id_838gat, id_827gat, id_781gat, id_712gat, id_527gat);
nand ( id_839gat, id_828gat, id_785gat, id_721gat, id_528gat);
not ( id_840gat, id_829gat);
nand ( id_841gat, id_815gat, id_593gat);
nor ( id_842gat, id_830gat, id_831gat);
nor ( id_843gat, id_832gat, id_833gat);
nor ( id_844gat, id_834gat, id_835gat);
nor ( id_845gat, id_334gat, id_836gat);
not ( id_846gat, id_837gat);
not ( id_847gat, id_838gat);
not ( id_848gat, id_839gat);
and ( id_849gat, id_735gat, id_841gat);
buf ( id_850gat, id_840gat);
and ( id_851gat, id_219gat, id_842gat);
and ( id_852gat, id_219gat, id_843gat);
and ( id_853gat, id_219gat, id_844gat);
nand ( id_854gat, id_845gat, id_772gat, id_696gat);
not ( id_855gat, id_846gat);
not ( id_856gat, id_847gat);
not ( id_857gat, id_848gat);
not ( id_858gat, id_849gat);
nor ( id_859gat, id_417gat, id_851gat);
nor ( id_860gat, id_332gat, id_852gat);
nor ( id_861gat, id_333gat, id_853gat);
not ( id_862gat, id_854gat);
buf ( id_863gat, id_855gat);
buf ( id_864gat, id_856gat);
buf ( id_865gat, id_857gat);
buf ( id_866gat, id_858gat);
nand ( id_867gat, id_859gat, id_769gat, id_669gat);
nand ( id_868gat, id_860gat, id_770gat, id_677gat);
nand ( id_869gat, id_861gat, id_771gat, id_686gat);
not ( id_870gat, id_862gat);
not ( id_871gat, id_867gat);
not ( id_872gat, id_868gat);
not ( id_873gat, id_869gat);
buf ( id_874gat, id_870gat);
not ( id_875gat, id_871gat);
not ( id_876gat, id_872gat);
not ( id_877gat, id_873gat);
buf ( id_878gat, id_875gat);
buf ( id_879gat, id_876gat);
buf ( id_880gat, id_877gat);

endmodule
