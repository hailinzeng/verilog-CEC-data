module c2670nr
( id_1 ,id_2 ,id_3 ,id_4 ,id_5 ,id_6 ,id_7 ,id_8 ,id_11 ,id_14 ,id_15 ,id_16 ,id_19 ,id_20 ,id_21 ,id_22 ,id_23 ,id_24 ,id_25 
,id_26 ,id_27 ,id_28 ,id_29 ,id_32 ,id_33 ,id_34 ,id_35 ,id_36 ,id_37 ,id_40 ,id_43 ,id_44 ,id_47 ,id_48 ,id_49 ,id_50 ,id_51 
,id_52 ,id_53 ,id_54 ,id_55 ,id_56 ,id_57 ,id_60 ,id_61 ,id_62 ,id_63 ,id_64 ,id_65 ,id_66 ,id_67 ,id_68 ,id_69 ,id_72 ,id_73 
,id_74 ,id_75 ,id_76 ,id_77 ,id_78 ,id_79 ,id_80 ,id_81 ,id_82 ,id_85 ,id_86 ,id_87 ,id_88 ,id_89 ,id_90 ,id_91 ,id_92 ,id_93 
,id_94 ,id_95 ,id_96 ,id_99 ,id_100 ,id_101 ,id_102 ,id_103 ,id_104 ,id_105 ,id_106 ,id_107 ,id_108 ,id_111 ,id_112 ,id_113 ,id_114 
,id_115 ,id_116 ,id_117 ,id_118 ,id_119 ,id_120 ,id_123 ,id_124 ,id_125 ,id_126 ,id_127 ,id_128 ,id_129 ,id_130 ,id_131 ,id_132 
,id_135 ,id_136 ,id_137 ,id_138 ,id_139 ,id_140 ,id_141 ,id_142 ,id_452 ,id_483 ,id_543 ,id_559 ,id_567 ,id_651 ,id_661 ,id_860 
,id_868 ,id_1083 ,id_1341 ,id_1348 ,id_1384 ,id_1956 ,id_1961 ,id_1966 ,id_1971 ,id_1976 ,id_1981 ,id_1986 ,id_1991 ,id_1996 
,id_2066 ,id_2067 ,id_2072 ,id_2078 ,id_2084 ,id_2090 ,id_2096 ,id_2100 ,id_2104 ,id_2105 ,id_2106 ,id_2427 ,id_2430 ,id_2435 
,id_2438 ,id_2443 ,id_2446 ,id_2451 ,id_2454 ,id_2474 ,id_2678 ,id_350 ,id_335 ,id_409 ,id_369 ,id_367 ,id_411 ,id_337 ,id_384 
,id_218 ,id_219 ,id_220 ,id_221 ,id_235 ,id_236 ,id_237 ,id_238 ,id_158 ,id_259 ,id_391 ,id_173 ,id_223 ,id_234 ,id_217 ,id_325 
,id_261 ,id_319 ,id_160 ,id_162 ,id_164 ,id_166 ,id_168 ,id_171 ,id_153 ,id_176 ,id_188 ,id_299 ,id_301 ,id_286 ,id_303 ,id_288 
,id_305 ,id_290 ,id_284 ,id_321 ,id_297 ,id_280 ,id_148 ,id_282 ,id_323 ,id_156 ,id_401 ,id_227 ,id_229 ,id_311 ,id_150 ,id_145 
,id_395 ,id_295 ,id_331 ,id_397 ,id_329 ,id_308 ,id_225 /*, id_231*/ );

input id_1, id_2, id_3, id_4, id_5, id_6, id_7, id_8, id_11, id_14, id_15, id_16, id_19, id_20, id_21, id_22, id_23, id_24, id_25, id_26, id_27, id_28, id_29, id_32, id_33, id_34, id_35, id_36, id_37, id_40, id_43, id_44, id_47, id_48, id_49, id_50, id_51, id_52, id_53, id_54, id_55, id_56, id_57, id_60, id_61, id_62, id_63, id_64, id_65, id_66, id_67, id_68, id_69, id_72, id_73, id_74, id_75, id_76, id_77, id_78, id_79, id_80, id_81, id_82, id_85, id_86, id_87, id_88, id_89, id_90, id_91, id_92, id_93, id_94, id_95, id_96, id_99, id_100, id_101, id_102, id_103, id_104, id_105, id_106, id_107, id_108, id_111, id_112, id_113, id_114, id_115, id_116, id_117, id_118, id_119, id_120, id_123, id_124, id_125, id_126, id_127, id_128, id_129, id_130, id_131, id_132, id_135, id_136, id_137, id_138, id_139, id_140, id_141, id_142, id_452, id_483, id_543, id_559, id_567, id_651, id_661, id_860, id_868, id_1083, id_1341, id_1348, id_1384, id_1956, id_1961, id_1966, id_1971, id_1976, id_1981, id_1986, id_1991, id_1996, id_2066, id_2067, id_2072, id_2078, id_2084, id_2090, id_2096, id_2100, id_2104, id_2105, id_2106, id_2427, id_2430, id_2435, id_2438, id_2443, id_2446, id_2451, id_2454, id_2474, id_2678;

output id_350, id_335, id_409, id_369, id_367, id_411, id_337, id_384, id_218, id_219, id_220, id_221, id_235, id_236, id_237, id_238, id_158, id_259, id_391, id_173, id_223, id_234, id_217, id_325, id_261, id_319, id_160, id_162, id_164, id_166, id_168, id_171, id_153, id_176, id_188, id_299, id_301, id_286, id_303, id_288, id_305, id_290, id_284, id_321, id_297, id_280, id_148, id_282, id_323, id_156, id_401, id_227, id_229, id_311, id_150, id_145, id_395, id_295, id_331, id_397, id_329, /*id_231,*/ id_308, id_225;

buf ( id_350, id_452);
buf ( id_335, id_452);
buf ( id_409, id_452);
and ( id_546, id_1, id_3);
not ( id_560, id_559);
buf ( id_369, id_1083);
buf ( id_367, id_1083);
not ( id_1385, id_1384);
buf ( id_411, id_2066);
buf ( id_337, id_2066);
buf ( id_384, id_2066);
and ( id_157, id_2090, id_2084, id_2078, id_2072);
not ( id_547, id_546);
not ( id_218, id_44);
not ( id_219, id_132);
not ( id_220, id_82);
not ( id_221, id_96);
not ( id_235, id_69);
not ( id_236, id_120);
not ( id_237, id_57);
not ( id_238, id_108);
and ( id_258, id_2, id_15, id_661);
buf ( id_480, id_661);
buf ( id_486, id_37);
buf ( id_654, id_452);
buf ( id_655, id_8);
buf ( id_658, id_8);
buf ( id_772, id_543);
buf ( id_795, id_651);
not ( id_865, id_860);
not ( id_875, id_868);
buf ( id_882, id_11);
and ( id_1251, id_132, id_82, id_96, id_44);
and ( id_1254, id_120, id_57, id_108, id_69);
buf ( id_1261, id_543);
buf ( id_1284, id_651);
not ( id_1344, id_1341);
not ( id_1351, id_1348);
buf ( id_1394, id_2104);
buf ( id_1418, id_2105);
not ( id_2433, id_2427);
not ( id_2434, id_2430);
not ( id_2441, id_2435);
not ( id_2442, id_2438);
not ( id_2449, id_2443);
not ( id_2450, id_2446);
not ( id_2478, id_2474);
buf ( id_1631, id_2104);
buf ( id_1655, id_2105);
buf ( id_1710, id_16);
buf ( id_1721, id_16);
not ( id_2682, id_2678);
and ( id_1955, id_7, id_661);
not ( id_1959, id_1956);
not ( id_1964, id_1961);
not ( id_1969, id_1966);
not ( id_1974, id_1971);
not ( id_1979, id_1976);
not ( id_1984, id_1981);
not ( id_1989, id_1986);
not ( id_1994, id_1991);
not ( id_1999, id_1996);
buf ( id_2001, id_29);
buf ( id_2012, id_29);
not ( id_2070, id_2067);
not ( id_2076, id_2072);
not ( id_2082, id_2078);
not ( id_2088, id_2084);
not ( id_2094, id_2090);
not ( id_2099, id_2096);
not ( id_2103, id_2100);
not ( id_2457, id_2451);
not ( id_2458, id_2454);
buf ( id_2461, id_1348);
buf ( id_2464, id_1341);
buf ( id_2471, id_1956);
buf ( id_2479, id_1966);
buf ( id_2482, id_1961);
buf ( id_2487, id_1976);
buf ( id_2490, id_1971);
buf ( id_2495, id_1986);
buf ( id_2498, id_1981);
buf ( id_2505, id_1996);
buf ( id_2508, id_1991);
buf ( id_2675, id_2067);
buf ( id_2683, id_2078);
buf ( id_2686, id_2072);
buf ( id_2691, id_2090);
buf ( id_2694, id_2084);
buf ( id_2699, id_2100);
buf ( id_2702, id_2096);
not ( id_158, id_157);
not ( id_259, id_258);
not ( id_487, id_486);
buf ( id_391, id_654);
nand ( id_1475, id_2430, id_2433);
nand ( id_1476, id_2427, id_2434);
nand ( id_1484, id_2438, id_2441);
nand ( id_1485, id_2435, id_2442);
nand ( id_1493, id_2446, id_2449);
nand ( id_1494, id_2443, id_2450);
nand ( id_2459, id_2454, id_2457);
nand ( id_2460, id_2451, id_2458);
and ( id_173, id_94, id_654);
and ( id_216, id_2106, id_1955);
not ( id_223, id_1955);
nand ( id_234, id_567, id_1955);
not ( id_1253, id_1251);
not ( id_1256, id_1254);
and ( id_558, id_1254, id_1251);
not ( id_784, id_772);
not ( id_807, id_795);
and ( id_821, id_80, id_772, id_795);
and ( id_825, id_68, id_772, id_795);
and ( id_829, id_79, id_772, id_795);
and ( id_833, id_78, id_772, id_795);
and ( id_837, id_77, id_772, id_795);
buf ( id_994, id_655);
not ( id_1273, id_1261);
not ( id_1296, id_1284);
and ( id_1310, id_76, id_1261, id_1284);
and ( id_1314, id_75, id_1261, id_1284);
and ( id_1318, id_74, id_1284);
and ( id_1322, id_73, id_1261, id_1284);
and ( id_1326, id_72, id_1261, id_1284);
not ( id_1406, id_1394);
not ( id_1430, id_1418);
and ( id_1444, id_114, id_1394, id_1418);
and ( id_1448, id_113, id_1394, id_1418);
and ( id_1452, id_112, id_1394, id_1418);
and ( id_1456, id_111, id_1394, id_1418);
nand ( id_1477, id_1475, id_1476);
nand ( id_1486, id_1484, id_1485);
nand ( id_1495, id_1493, id_1494);
not ( id_2477, id_2471);
nand ( id_1499, id_2471, id_2478);
not ( id_2485, id_2479);
not ( id_2486, id_2482);
not ( id_2493, id_2487);
not ( id_2494, id_2490);
not ( id_1643, id_1631);
not ( id_1667, id_1655);
and ( id_1681, id_118, id_1631, id_1655);
and ( id_1685, id_107, id_1631, id_1655);
and ( id_1689, id_117, id_1631, id_1655);
and ( id_1693, id_116, id_1631, id_1655);
and ( id_1697, id_115, id_1631, id_1655);
not ( id_1716, id_1710);
not ( id_1728, id_1721);
not ( id_2681, id_2675);
nand ( id_1776, id_2675, id_2682);
not ( id_2689, id_2683);
not ( id_2690, id_2686);
not ( id_2697, id_2691);
not ( id_2698, id_2694);
buf ( id_1893, id_658);
not ( id_2007, id_2001);
not ( id_2018, id_2012);
not ( id_2467, id_2461);
not ( id_2468, id_2464);
not ( id_2501, id_2495);
not ( id_2502, id_2498);
not ( id_2511, id_2505);
not ( id_2512, id_2508);
nand ( id_2518, id_2459, id_2460);
buf ( id_2551, id_1344);
buf ( id_2559, id_1351);
buf ( id_2567, id_1959);
buf ( id_2575, id_1964);
buf ( id_2583, id_1969);
buf ( id_2591, id_1974);
buf ( id_2599, id_1979);
buf ( id_2607, id_1984);
buf ( id_2615, id_1989);
buf ( id_2623, id_1994);
not ( id_2705, id_2699);
not ( id_2706, id_2702);
buf ( id_2735, id_1999);
buf ( id_2743, id_2070);
buf ( id_2751, id_2076);
buf ( id_2759, id_2082);
buf ( id_2767, id_2088);
buf ( id_2775, id_2094);
not ( id_217, id_216);
and ( id_550, id_2106, id_1253);
and ( id_552, id_567, id_1256);
buf ( id_325, id_558);
buf ( id_894, id_882);
nand ( id_1498, id_2474, id_2477);
nand ( id_1507, id_2482, id_2485);
nand ( id_1508, id_2479, id_2486);
nand ( id_1516, id_2490, id_2493);
nand ( id_1517, id_2487, id_2494);
nand ( id_1775, id_2678, id_2681);
nand ( id_1784, id_2686, id_2689);
nand ( id_1785, id_2683, id_2690);
nand ( id_1793, id_2694, id_2697);
nand ( id_1794, id_2691, id_2698);
nand ( id_2469, id_2464, id_2467);
nand ( id_2470, id_2461, id_2468);
nand ( id_2503, id_2498, id_2501);
nand ( id_2504, id_2495, id_2502);
nand ( id_2513, id_2508, id_2511);
nand ( id_2514, id_2505, id_2512);
nand ( id_2707, id_2702, id_2705);
nand ( id_2708, id_2699, id_2706);
not ( id_261, id_558);
not ( id_551, id_550);
not ( id_553, id_552);
and ( id_818, id_93, id_784, id_807);
and ( id_819, id_55, id_772, id_807);
and ( id_820, id_67, id_784, id_795);
and ( id_822, id_81, id_784, id_807);
and ( id_823, id_43, id_772, id_807);
and ( id_824, id_56, id_784, id_795);
and ( id_826, id_92, id_784, id_807);
and ( id_827, id_54, id_772, id_807);
and ( id_828, id_66, id_784, id_795);
and ( id_830, id_91, id_784, id_807);
and ( id_831, id_53, id_772, id_807);
and ( id_832, id_65, id_784, id_795);
and ( id_834, id_90, id_784, id_807);
and ( id_835, id_52, id_772, id_807);
and ( id_836, id_64, id_784, id_795);
and ( id_1307, id_89, id_1273, id_1296);
and ( id_1308, id_51, id_1261, id_1296);
and ( id_1309, id_63, id_1273, id_1284);
and ( id_1311, id_88, id_1273, id_1296);
and ( id_1312, id_50, id_1261, id_1296);
and ( id_1313, id_62, id_1273, id_1284);
and ( id_1315, id_87, id_1273);
and ( id_1316, id_49, id_1261, id_1296);
and ( id_1317, id_1273, id_1284);
and ( id_1319, id_86, id_1273, id_1296);
and ( id_1320, id_48, id_1261, id_1296);
and ( id_1321, id_61, id_1273, id_1284);
and ( id_1323, id_85, id_1273, id_1296);
and ( id_1324, id_47, id_1261, id_1296);
and ( id_1325, id_60, id_1273, id_1284);
and ( id_1441, id_138, id_1406, id_1430);
and ( id_1442, id_102, id_1394, id_1430);
and ( id_1443, id_126, id_1406, id_1418);
and ( id_1445, id_137, id_1406, id_1430);
and ( id_1446, id_101, id_1394, id_1430);
and ( id_1447, id_125, id_1406, id_1418);
and ( id_1449, id_136, id_1406, id_1430);
and ( id_1450, id_100, id_1394, id_1430);
and ( id_1451, id_124, id_1406, id_1418);
and ( id_1453, id_135, id_1406, id_1430);
and ( id_1454, id_99, id_1394, id_1430);
and ( id_1455, id_123, id_1406, id_1418);
not ( id_1481, id_1477);
not ( id_1490, id_1486);
nand ( id_1500, id_1498, id_1499);
nand ( id_1509, id_1507, id_1508);
nand ( id_1518, id_1516, id_1517);
buf ( id_1521, id_1495);
buf ( id_1525, id_1495);
not ( id_2557, id_2551);
not ( id_2565, id_2559);
not ( id_2573, id_2567);
not ( id_2581, id_2575);
not ( id_2589, id_2583);
not ( id_2597, id_2591);
not ( id_2605, id_2599);
not ( id_2613, id_2607);
not ( id_2621, id_2615);
not ( id_2629, id_2623);
and ( id_1678, id_142, id_1643, id_1667);
and ( id_1679, id_106, id_1631, id_1667);
and ( id_1680, id_130, id_1643, id_1655);
and ( id_1682, id_131, id_1643, id_1667);
and ( id_1683, id_95, id_1631, id_1667);
and ( id_1684, id_119, id_1643, id_1655);
and ( id_1686, id_141, id_1643, id_1667);
and ( id_1687, id_105, id_1631, id_1667);
and ( id_1688, id_129, id_1643, id_1655);
and ( id_1690, id_140, id_1643, id_1667);
and ( id_1691, id_104, id_1631, id_1667);
and ( id_1692, id_128, id_1643, id_1655);
and ( id_1694, id_139, id_1643, id_1667);
and ( id_1695, id_103, id_1631, id_1667);
and ( id_1696, id_127, id_1643, id_1655);
and ( id_1734, id_19, id_1716);
and ( id_1736, id_4, id_1716);
and ( id_1738, id_20, id_1716);
and ( id_1740, id_5, id_1716);
and ( id_1742, id_21, id_1728);
and ( id_1744, id_22, id_1728);
and ( id_1746, id_23, id_1728);
and ( id_1748, id_6, id_1728);
and ( id_1750, id_24, id_1728);
nand ( id_1777, id_1775, id_1776);
nand ( id_1786, id_1784, id_1785);
nand ( id_1795, id_1793, id_1794);
and ( id_2023, id_25, id_2007);
and ( id_2025, id_32, id_2007);
and ( id_2027, id_26, id_2007);
and ( id_2029, id_33, id_2007);
and ( id_2031, id_27, id_2018);
and ( id_2033, id_34, id_2018);
and ( id_2035, id_35, id_2018);
and ( id_2037, id_28, id_2018);
not ( id_2741, id_2735);
not ( id_2749, id_2743);
not ( id_2757, id_2751);
not ( id_2765, id_2759);
not ( id_2773, id_2767);
not ( id_2781, id_2775);
nand ( id_2515, id_2469, id_2470);
not ( id_2522, id_2518);
nand ( id_2525, id_2513, id_2514);
nand ( id_2528, id_2503, id_2504);
nand ( id_2730, id_2707, id_2708);
and ( id_554, id_551, id_553);
or ( id_838, id_818, id_819, id_820, id_821);
or ( id_841, id_822, id_823, id_824, id_825);
or ( id_846, id_826, id_827, id_828, id_829);
or ( id_854, id_830, id_831, id_832, id_833);
or ( id_857, id_834, id_835, id_836, id_837);
or ( id_1327, id_1307, id_1308, id_1309, id_1310);
or ( id_1329, id_1311, id_1312, id_1313, id_1314);
or ( id_1331, id_1315, id_1316, id_1317, id_1318);
or ( id_1333, id_1319, id_1320, id_1321, id_1322);
or ( id_1335, id_1323, id_1324, id_1325, id_1326);
or ( id_1461, id_1441, id_1442, id_1443, id_1444);
or ( id_1464, id_1445, id_1446, id_1447, id_1448);
or ( id_1467, id_1449, id_1450, id_1451, id_1452);
or ( id_1470, id_1453, id_1454, id_1455, id_1456);
or ( id_1698, id_1682, id_1683, id_1684, id_1685);
or ( id_1701, id_1686, id_1687, id_1688, id_1689);
or ( id_1704, id_1690, id_1691, id_1692, id_1693);
or ( id_1707, id_1694, id_1695, id_1696, id_1697);
or ( id_2634, id_1678, id_1679, id_1680, id_1681);
buf ( id_319, id_554);
not ( id_1504, id_1500);
not ( id_1513, id_1509);
not ( id_1524, id_1521);
not ( id_1528, id_1525);
buf ( id_1529, id_1518);
buf ( id_1533, id_1518);
and ( id_1538, id_1486, id_1477, id_1521);
and ( id_1541, id_1490, id_1481, id_1525);
not ( id_1781, id_1777);
not ( id_1790, id_1786);
buf ( id_1806, id_1795);
buf ( id_1810, id_1795);
not ( id_2734, id_2730);
not ( id_2521, id_2515);
nand ( id_2524, id_2515, id_2522);
not ( id_2531, id_2525);
not ( id_2532, id_2528);
and ( id_144, id_838, id_860);
buf ( id_147, id_846);
buf ( id_152, id_841);
not ( id_160, id_1464);
not ( id_162, id_1467);
not ( id_164, id_1461);
not ( id_166, id_1329);
not ( id_168, id_1327);
not ( id_171, id_857);
and ( id_175, id_480, id_483, id_36, id_554);
and ( id_187, id_480, id_483, id_554, id_547);
buf ( id_516, id_838);
not ( id_852, id_846);
and ( id_885, id_841, id_875);
and ( id_887, id_846, id_875);
and ( id_893, id_1327, id_868);
not ( id_1028, id_838);
not ( id_1031, id_841);
not ( id_1035, id_846);
buf ( id_1041, id_854);
buf ( id_1049, id_857);
buf ( id_1057, id_1327);
buf ( id_1060, id_1329);
buf ( id_1066, id_1331);
buf ( id_1072, id_1333);
buf ( id_1078, id_1335);
nand ( id_1213, id_2099, id_1470);
not ( id_1218, id_2103);
buf ( id_1250, id_1704);
and ( id_1387, id_1461, id_1385);
not ( id_1389, id_1464);
and ( id_1537, id_1481, id_1486, id_1524);
and ( id_1540, id_1477, id_1490, id_1528);
and ( id_1735, id_841, id_1710);
and ( id_1737, id_846, id_1710);
and ( id_1739, id_854, id_1710);
and ( id_1741, id_857, id_1710);
and ( id_1743, id_1327, id_1721);
and ( id_1745, id_1329, id_1721);
and ( id_1747, id_1331, id_1721);
and ( id_1749, id_1333, id_1721);
and ( id_1751, id_1335, id_1721);
not ( id_2638, id_2634);
and ( id_2024, id_1698, id_2001);
and ( id_2026, id_1701, id_2001);
and ( id_2028, id_1704, id_2001);
and ( id_2030, id_1707, id_2001);
and ( id_2032, id_1461, id_2012);
and ( id_2034, id_1464, id_2012);
and ( id_2036, id_1467, id_2012);
and ( id_2038, id_1470, id_2012);
buf ( id_2154, id_841);
nand ( id_2523, id_2518, id_2521);
nand ( id_2533, id_2528, id_2531);
nand ( id_2534, id_2525, id_2532);
buf ( id_2631, id_1698);
buf ( id_2639, id_1704);
buf ( id_2642, id_1701);
buf ( id_2647, id_1461);
buf ( id_2650, id_1707);
buf ( id_2655, id_1467);
buf ( id_2658, id_1464);
buf ( id_2668, id_1470);
or ( id_153, id_865, id_152);
not ( id_176, id_175);
not ( id_188, id_187);
buf ( id_299, id_1041);
buf ( id_301, id_1049);
buf ( id_286, id_1057);
buf ( id_303, id_1060);
buf ( id_288, id_1066);
buf ( id_305, id_1072);
buf ( id_290, id_1078);
not ( id_1532, id_1529);
not ( id_1536, id_1533);
nor ( id_1539, id_1537, id_1538);
nor ( id_1542, id_1540, id_1541);
and ( id_1544, id_1509, id_1500, id_1529);
and ( id_1547, id_1513, id_1504, id_1533);
or ( id_2065, id_2037, id_2038);
not ( id_1809, id_1806);
not ( id_1813, id_1810);
and ( id_1821, id_1786, id_1777, id_1806);
and ( id_1824, id_1790, id_1781, id_1810);
nand ( id_2538, id_2523, id_2524);
nand ( id_2546, id_2533, id_2534);
or ( id_2554, id_1734, id_1735);
or ( id_2562, id_1736, id_1737);
or ( id_2570, id_1738, id_1739);
or ( id_2578, id_1740, id_1741);
or ( id_2586, id_1742, id_1743);
or ( id_2594, id_1744, id_1745);
or ( id_2602, id_1746, id_1747);
or ( id_2610, id_1748, id_1749);
or ( id_2618, id_1750, id_1751);
or ( id_2626, id_2023, id_2024);
or ( id_2738, id_2025, id_2026);
or ( id_2746, id_2027, id_2028);
or ( id_2754, id_2029, id_2030);
or ( id_2762, id_2031, id_2032);
or ( id_2770, id_2033, id_2034);
or ( id_2778, id_2035, id_2036);
and ( id_456, id_1389, id_1387, id_40);
nand ( id_562, id_560, id_852);
and ( id_883, id_516, id_875);
and ( id_889, id_1049, id_868);
and ( id_891, id_1041, id_875);
not ( id_1043, id_1041);
not ( id_1051, id_1049);
not ( id_1062, id_1060);
not ( id_1068, id_1066);
not ( id_1074, id_1072);
not ( id_1080, id_1078);
and ( id_1225, id_2099, id_1213);
and ( id_1227, id_1213, id_1470);
buf ( id_1234, id_1218);
and ( id_1543, id_1504, id_1509, id_1532);
and ( id_1546, id_1500, id_1513, id_1536);
not ( id_2637, id_2631);
nand ( id_1753, id_2631, id_2638);
not ( id_2645, id_2639);
not ( id_2646, id_2642);
not ( id_2653, id_2647);
not ( id_2654, id_2650);
and ( id_1820, id_1781, id_1786, id_1809);
and ( id_1823, id_1777, id_1790, id_1813);
buf ( id_2107, id_1031);
buf ( id_2110, id_1028);
buf ( id_2118, id_1035);
not ( id_2123, id_1057);
not ( id_2151, id_852);
not ( id_2158, id_2154);
buf ( id_2161, id_1031);
buf ( id_2164, id_1028);
buf ( id_2172, id_1035);
buf ( id_2235, id_516);
buf ( id_2350, id_1035);
nand ( id_2535, id_1542, id_1539);
not ( id_2661, id_2655);
not ( id_2662, id_2658);
not ( id_2672, id_2668);
and ( id_468, id_40, id_1389);
or ( id_897, id_887, id_889);
or ( id_898, id_891, id_893);
or ( id_1228, id_1225, id_1227);
buf ( id_1235, id_1234);
nor ( id_1545, id_1543, id_1544);
nor ( id_1548, id_1546, id_1547);
not ( id_2542, id_2538);
not ( id_2550, id_2546);
nand ( id_1561, id_2554, id_2557);
not ( id_2558, id_2554);
nand ( id_1565, id_2562, id_2565);
not ( id_2566, id_2562);
nand ( id_1569, id_2570, id_2573);
not ( id_2574, id_2570);
nand ( id_1573, id_2578, id_2581);
not ( id_2582, id_2578);
nand ( id_1577, id_2586, id_2589);
not ( id_2590, id_2586);
nand ( id_1581, id_2594, id_2597);
not ( id_2598, id_2594);
nand ( id_1585, id_2602, id_2605);
not ( id_2606, id_2602);
nand ( id_1589, id_2610, id_2613);
not ( id_2614, id_2610);
nand ( id_1593, id_2618, id_2621);
not ( id_2622, id_2618);
nand ( id_1597, id_2626, id_2629);
not ( id_2630, id_2626);
nand ( id_1752, id_2634, id_2637);
nand ( id_1761, id_2642, id_2645);
nand ( id_1762, id_2639, id_2646);
nand ( id_1770, id_2650, id_2653);
nand ( id_1771, id_2647, id_2654);
nor ( id_1822, id_1820, id_1821);
nor ( id_1825, id_1823, id_1824);
nand ( id_2039, id_2738, id_2741);
not ( id_2742, id_2738);
nand ( id_2043, id_2746, id_2749);
not ( id_2750, id_2746);
nand ( id_2047, id_2754, id_2757);
not ( id_2758, id_2754);
nand ( id_2051, id_2762, id_2765);
not ( id_2766, id_2762);
nand ( id_2055, id_2770, id_2773);
not ( id_2774, id_2770);
nand ( id_2059, id_2778, id_2781);
not ( id_2782, id_2778);
nand ( id_2663, id_2658, id_2661);
nand ( id_2664, id_2655, id_2662);
not ( id_2674, id_2672);
and ( id_146, id_562, id_865);
not ( id_462, id_456);
not ( id_2113, id_2107);
not ( id_2114, id_2110);
not ( id_2122, id_2118);
not ( id_2129, id_2123);
buf ( id_592, id_562);
not ( id_2167, id_2161);
not ( id_2168, id_2164);
not ( id_2176, id_2172);
not ( id_2241, id_2235);
and ( id_886, id_562, id_868);
buf ( id_284, id_897);
buf ( id_321, id_897);
buf ( id_297, id_898);
buf ( id_280, id_898);
buf ( id_995, id_456);
not ( id_1006, id_456);
nand ( id_1550, id_2535, id_2542);
not ( id_2541, id_2535);
nand ( id_1562, id_2551, id_2558);
nand ( id_1566, id_2559, id_2566);
nand ( id_1570, id_2567, id_2574);
nand ( id_1574, id_2575, id_2582);
nand ( id_1578, id_2583, id_2590);
nand ( id_1582, id_2591, id_2598);
nand ( id_1586, id_2599, id_2606);
nand ( id_1590, id_2607, id_2614);
nand ( id_1594, id_2615, id_2622);
nand ( id_1598, id_2623, id_2630);
nand ( id_1754, id_1752, id_1753);
nand ( id_1763, id_1761, id_1762);
nand ( id_1772, id_1770, id_1771);
nand ( id_2040, id_2735, id_2742);
nand ( id_2044, id_2743, id_2750);
nand ( id_2048, id_2751, id_2758);
nand ( id_2052, id_2759, id_2766);
nand ( id_2056, id_2767, id_2774);
nand ( id_2060, id_2775, id_2782);
buf ( id_2115, id_1043);
buf ( id_2126, id_1051);
buf ( id_2131, id_1068);
buf ( id_2134, id_1062);
buf ( id_2141, id_1080);
buf ( id_2144, id_1074);
not ( id_2157, id_2151);
nand ( id_2160, id_2151, id_2158);
buf ( id_2169, id_1043);
buf ( id_2177, id_1068);
buf ( id_2180, id_1062);
buf ( id_2187, id_1080);
buf ( id_2190, id_1074);
not ( id_2207, id_562);
buf ( id_2342, id_1043);
buf ( id_2422, id_1051);
nand ( id_2543, id_1548, id_1545);
not ( id_2709, id_2674);
nand ( id_2712, id_2663, id_2664);
nand ( id_2727, id_1825, id_1822);
or ( id_148, id_146, id_147);
nand ( id_569, id_2110, id_2113);
nand ( id_570, id_2107, id_2114);
nand ( id_599, id_2164, id_2167);
nand ( id_600, id_2161, id_2168);
or ( id_896, id_885, id_886);
nand ( id_1549, id_2538, id_2541);
not ( id_1243, id_1228);
not ( id_1245, id_1235);
buf ( id_1257, id_468);
buf ( id_1258, id_468);
nand ( id_1563, id_1561, id_1562);
nand ( id_1567, id_1565, id_1566);
nand ( id_1571, id_1569, id_1570);
nand ( id_1575, id_1573, id_1574);
nand ( id_1579, id_1577, id_1578);
nand ( id_1583, id_1581, id_1582);
nand ( id_1587, id_1585, id_1586);
nand ( id_1591, id_1589, id_1590);
nand ( id_1595, id_1593, id_1594);
nand ( id_1599, id_1597, id_1598);
nand ( id_2041, id_2039, id_2040);
nand ( id_2045, id_2043, id_2044);
nand ( id_2049, id_2047, id_2048);
nand ( id_2053, id_2051, id_2052);
nand ( id_2057, id_2055, id_2056);
nand ( id_2061, id_2059, id_2060);
nand ( id_2159, id_2154, id_2157);
nand ( id_571, id_569, id_570);
not ( id_2121, id_2115);
nand ( id_579, id_2115, id_2122);
nand ( id_587, id_2126, id_2129);
not ( id_2130, id_2126);
not ( id_596, id_592);
nand ( id_601, id_599, id_600);
not ( id_2175, id_2169);
nand ( id_609, id_2169, id_2176);
buf ( id_1014, id_1057);
buf ( id_1018, id_1060);
and ( id_717, id_1078, id_1006);
and ( id_723, id_1698, id_1006);
and ( id_729, id_1701, id_1006);
and ( id_735, id_1250, id_1006);
buf ( id_282, id_896);
buf ( id_323, id_896);
not ( id_999, id_995);
nand ( id_1091, id_1549, id_1550);
buf ( id_1337, id_462);
not ( id_2549, id_2543);
nand ( id_1552, id_2543, id_2550);
not ( id_1600, id_1599);
not ( id_1596, id_1595);
not ( id_1592, id_1591);
not ( id_1588, id_1587);
not ( id_1584, id_1583);
not ( id_1580, id_1579);
not ( id_1576, id_1575);
not ( id_1572, id_1571);
not ( id_1568, id_1567);
not ( id_1564, id_1563);
not ( id_2062, id_2061);
not ( id_2058, id_2057);
not ( id_2054, id_2053);
not ( id_2050, id_2049);
not ( id_2046, id_2045);
not ( id_2042, id_2041);
not ( id_1758, id_1754);
not ( id_1767, id_1763);
buf ( id_1798, id_1772);
buf ( id_1802, id_1772);
not ( id_2733, id_2727);
nand ( id_1829, id_2727, id_2734);
not ( id_2137, id_2131);
not ( id_2138, id_2134);
not ( id_2147, id_2141);
not ( id_2148, id_2144);
not ( id_2183, id_2177);
not ( id_2184, id_2180);
not ( id_2193, id_2187);
not ( id_2194, id_2190);
nand ( id_2210, id_2159, id_2160);
not ( id_2213, id_2207);
not ( id_2715, id_2709);
not ( id_2716, id_2712);
nand ( id_578, id_2118, id_2121);
nand ( id_588, id_2123, id_2130);
nand ( id_608, id_2172, id_2175);
buf ( id_1005, id_1257);
not ( id_1092, id_1091);
nand ( id_1551, id_2546, id_2549);
and ( id_1554, id_1600, id_1596, id_1592, id_1588, id_1584);
and ( id_1555, id_1580, id_1576, id_1572, id_1568, id_1564);
and ( id_1557, id_2065, id_2062);
and ( id_1558, id_2058, id_2054, id_2050, id_2046, id_2042);
nand ( id_1828, id_2730, id_2733);
buf ( id_1907, id_1258);
nand ( id_2139, id_2134, id_2137);
nand ( id_2140, id_2131, id_2138);
nand ( id_2149, id_2144, id_2147);
nand ( id_2150, id_2141, id_2148);
nand ( id_2185, id_2180, id_2183);
nand ( id_2186, id_2177, id_2184);
nand ( id_2195, id_2190, id_2193);
nand ( id_2196, id_2187, id_2194);
nand ( id_2717, id_2712, id_2715);
nand ( id_2718, id_2709, id_2716);
buf ( id_154, id_1245);
buf ( id_155, id_1243);
not ( id_575, id_571);
nand ( id_580, id_578, id_579);
nand ( id_589, id_587, id_588);
not ( id_605, id_601);
nand ( id_610, id_608, id_609);
and ( id_705, id_1066, id_999);
and ( id_711, id_1072, id_999);
and ( id_1093, id_1092, id_14);
nand ( id_1553, id_1551, id_1552);
and ( id_1556, id_1554, id_1555);
and ( id_1559, id_1557, id_1558);
buf ( id_1601, id_1337);
not ( id_1801, id_1798);
not ( id_1805, id_1802);
and ( id_1815, id_1763, id_1754, id_1798);
and ( id_1818, id_1767, id_1758, id_1802);
nand ( id_1830, id_1828, id_1829);
buf ( id_1898, id_1337);
buf ( id_1912, id_1337);
nand ( id_2197, id_2149, id_2150);
nand ( id_2200, id_2139, id_2140);
not ( id_2214, id_2210);
nand ( id_2215, id_2210, id_2213);
nand ( id_2217, id_2195, id_2196);
nand ( id_2220, id_2185, id_2186);
nand ( id_2722, id_2717, id_2718);
nand ( id_156, id_154, id_155);
buf ( id_693, id_1014);
buf ( id_699, id_1018);
and ( id_707, id_705, id_994);
and ( id_713, id_711, id_994);
and ( id_719, id_717, id_1005);
and ( id_725, id_723, id_1005);
and ( id_731, id_729, id_1005);
and ( id_737, id_735, id_1005);
buf ( id_401, id_1093);
and ( id_1560, id_1556, id_1559, id_894);
and ( id_1814, id_1758, id_1763, id_1801);
and ( id_1817, id_1754, id_1767, id_1805);
nand ( id_2216, id_2207, id_2214);
not ( id_227, id_1830);
not ( id_229, id_1553);
not ( id_584, id_580);
buf ( id_613, id_589);
buf ( id_617, id_589);
buf ( id_621, id_610);
buf ( id_625, id_610);
and ( id_695, id_693, id_994);
and ( id_701, id_699, id_994);
not ( id_708, id_707);
not ( id_714, id_713);
not ( id_720, id_719);
not ( id_726, id_725);
not ( id_732, id_731);
not ( id_738, id_737);
not ( id_1087, id_1093);
and ( id_1108, id_1344, id_1601);
buf ( id_311, id_1560);
not ( id_1607, id_1601);
and ( id_1615, id_1351, id_1601);
and ( id_1619, id_1959, id_1601);
and ( id_1623, id_1964, id_1601);
nor ( id_1816, id_1814, id_1815);
nor ( id_1819, id_1817, id_1818);
not ( id_2726, id_2722);
not ( id_1904, id_1898);
and ( id_1920, id_1969, id_1898);
and ( id_1925, id_1974, id_1898);
and ( id_1928, id_1979, id_1898);
and ( id_1930, id_1984, id_1898);
and ( id_1932, id_1989, id_1912);
and ( id_1934, id_1994, id_1912);
and ( id_1936, id_1999, id_1912);
and ( id_1938, id_2070, id_1912);
not ( id_2203, id_2197);
not ( id_2204, id_2200);
not ( id_2223, id_2217);
not ( id_2224, id_2220);
nand ( id_2238, id_2215, id_2216);
not ( id_150, id_1560);
not ( id_696, id_695);
not ( id_702, id_701);
and ( id_1943, id_1928, id_1893);
and ( id_1945, id_1930, id_1893);
and ( id_1947, id_1932, id_1907);
and ( id_1949, id_1934, id_1907);
and ( id_1951, id_1936, id_1907);
and ( id_1953, id_1938, id_1907);
nand ( id_2205, id_2200, id_2203);
nand ( id_2206, id_2197, id_2204);
nand ( id_2225, id_2220, id_2223);
nand ( id_2226, id_2217, id_2224);
nand ( id_2719, id_1819, id_1816);
not ( id_616, id_613);
not ( id_620, id_617);
not ( id_624, id_621);
not ( id_628, id_625);
and ( id_630, id_580, id_571, id_613);
and ( id_633, id_584, id_575, id_617);
and ( id_636, id_601, id_592, id_621);
and ( id_639, id_605, id_596, id_625);
nand ( id_645, id_2238, id_2241);
not ( id_2242, id_2238);
and ( id_1107, id_1999, id_1607);
and ( id_1614, id_2070, id_1607);
and ( id_1617, id_2076, id_1607);
and ( id_1621, id_2082, id_1607);
and ( id_1918, id_2088, id_1904);
and ( id_1923, id_2094, id_1904);
nand ( id_2230, id_2205, id_2206);
nand ( id_2246, id_2225, id_2226);
buf ( id_2358, id_738);
buf ( id_2366, id_732);
buf ( id_2374, id_726);
buf ( id_2382, id_720);
buf ( id_2390, id_714);
buf ( id_2398, id_708);
and ( id_629, id_575, id_580, id_616);
and ( id_632, id_571, id_584, id_620);
and ( id_635, id_596, id_601, id_624);
and ( id_638, id_592, id_605, id_628);
nand ( id_646, id_2235, id_2242);
nand ( id_1827, id_2719, id_2726);
or ( id_1109, id_1107, id_1108);
and ( id_1125, id_1953, id_738);
and ( id_1133, id_1951, id_732);
and ( id_1140, id_1949, id_726);
and ( id_1142, id_720, id_1947);
and ( id_1155, id_1945, id_714);
and ( id_1164, id_1943, id_708);
or ( id_1624, id_1614, id_1615);
or ( id_1626, id_1617, id_1619);
or ( id_1628, id_1621, id_1623);
not ( id_2725, id_2719);
or ( id_1921, id_1918, id_1920);
or ( id_1926, id_1923, id_1925);
buf ( id_2355, id_1953);
buf ( id_2363, id_1951);
buf ( id_2371, id_1949);
buf ( id_2379, id_1947);
buf ( id_2387, id_1945);
buf ( id_2395, id_1943);
buf ( id_2406, id_702);
buf ( id_2414, id_696);
nand ( id_647, id_645, id_646);
nor ( id_631, id_629, id_630);
nor ( id_634, id_632, id_633);
nor ( id_637, id_635, id_636);
nor ( id_640, id_638, id_639);
not ( id_2234, id_2230);
not ( id_2250, id_2246);
nand ( id_1826, id_2722, id_2725);
and ( id_1110, id_1109, id_1031);
and ( id_1939, id_1921, id_1893);
and ( id_1941, id_1926, id_1893);
and ( id_143, id_647, id_865);
nand ( id_686, id_1826, id_1827);
and ( id_1104, id_1626, id_1043);
and ( id_1106, id_1624, id_1035);
not ( id_1118, id_2355);
not ( id_1127, id_2363);
not ( id_1135, id_2371);
not ( id_1144, id_2379);
not ( id_1147, id_2387);
not ( id_1157, id_2395);
and ( id_1184, id_1628, id_1051);
nand ( id_2227, id_634, id_631);
nand ( id_2243, id_640, id_637);
buf ( id_2339, id_1626);
buf ( id_2347, id_1624);
buf ( id_2419, id_1628);
or ( id_145, id_143, id_144);
not ( id_687, id_686);
not ( id_1117, id_2358);
not ( id_1126, id_2366);
not ( id_1134, id_2374);
not ( id_1143, id_2382);
not ( id_1146, id_2390);
not ( id_1156, id_2398);
and ( id_1172, id_1941, id_702);
and ( id_1179, id_1939, id_696);
buf ( id_2403, id_1941);
buf ( id_2411, id_1939);
not ( id_2233, id_2227);
nand ( id_642, id_2227, id_2234);
not ( id_2249, id_2243);
nand ( id_649, id_2243, id_2250);
and ( id_688, id_687, id_487);
not ( id_1099, id_2339);
not ( id_1115, id_2347);
nand ( id_1119, id_1117, id_1118);
nand ( id_1128, id_1126, id_1127);
nand ( id_1136, id_1134, id_1135);
nand ( id_1145, id_1143, id_1144);
nand ( id_1148, id_1146, id_1147);
nand ( id_1158, id_1156, id_1157);
not ( id_1181, id_2419);
nand ( id_641, id_2230, id_2233);
nand ( id_648, id_2246, id_2249);
buf ( id_395, id_688);
not ( id_1098, id_2342);
not ( id_1114, id_2350);
not ( id_1166, id_2403);
not ( id_1174, id_2411);
not ( id_1180, id_2422);
nand ( id_643, id_641, id_642);
nand ( id_650, id_648, id_649);
not ( id_690, id_688);
nand ( id_1100, id_1098, id_1099);
nand ( id_1112, id_1114, id_1115);
not ( id_1165, id_2406);
not ( id_1173, id_2414);
nand ( id_1182, id_1180, id_1181);
and ( id_1185, id_1128, id_1145, id_1136, id_1119);
and ( id_1187, id_1119, id_1133);
and ( id_1188, id_1128, id_1119, id_1140);
and ( id_1189, id_1136, id_1119, id_1142, id_1128);
and ( id_1195, id_1148, id_1164);
and ( id_1196, id_1158, id_1148, id_1172);
not ( id_644, id_643);
and ( id_884, id_650, id_868);
nand ( id_1167, id_1165, id_1166);
nand ( id_1175, id_1173, id_1174);
not ( id_1186, id_1185);
or ( id_1190, id_1125, id_1187, id_1188, id_1189);
or ( id_895, id_883, id_884);
and ( id_1025, id_644, id_487);
and ( id_1111, id_1100, id_1106);
and ( id_1113, id_1112, id_1100, id_1110);
buf ( id_295, id_895);
buf ( id_331, id_895);
buf ( id_397, id_1025);
or ( id_1116, id_1104, id_1111, id_1113);
and ( id_1194, id_1158, id_1182, id_1167, id_1148, id_1175);
and ( id_1197, id_1167, id_1148, id_1179, id_1158);
and ( id_1198, id_1175, id_1167, id_1148, id_1184, id_1158);
not ( id_1027, id_1025);
or ( id_1199, id_1155, id_1195, id_1196, id_1197, id_1198);
and ( id_1200, id_1194, id_1116);
not ( id_1205, id_1186);
and ( id_1085, id_690, id_1027, id_1830);
or ( id_1201, id_1199, id_1200);
and ( id_1207, id_1205, id_1201);
buf ( id_1206, id_1190);
or ( id_1208, id_1206, id_1207);
buf ( id_329, id_1208);
// ( id_231, ???);//
and ( id_1088, id_1553, id_1087);
and ( id_1089, id_1085, id_1088, id_554);
buf ( id_308, id_1089);
not ( id_225, id_1089);

endmodule
