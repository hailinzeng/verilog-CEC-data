module c7552nr
( id_1 ,id_5 ,id_9 ,id_12 ,id_15 ,id_18 ,id_23 ,id_26 ,id_29 ,id_32 ,id_35 ,id_38 ,id_41 ,id_44 ,id_47 ,id_50 ,id_53 ,id_54 ,id_55 ,id_56 ,id_57 ,id_58 ,id_59 ,id_60 ,id_61 ,id_62 ,id_63 ,id_64 ,id_65 ,id_66 ,id_69 ,id_70 ,id_73 ,id_74 ,id_75 ,id_76 ,id_77 ,id_78 ,id_79 ,id_80 ,id_81 ,id_82 ,id_83 ,id_84 ,id_85 ,id_86 ,id_87 ,id_88 ,id_89 ,id_94 ,id_97 ,id_100 ,id_103 ,id_106 ,id_109 ,id_110 ,id_111 ,id_112 ,id_113 ,id_114 ,id_115 ,id_118 ,id_121 ,id_124 ,id_127 ,id_130 ,id_133 ,id_134 ,id_135 ,id_138 ,id_141 ,id_144 ,id_147 ,id_150 ,id_151 ,id_152 ,id_153 ,id_154 ,id_155 ,id_156 ,id_157 ,id_158 ,id_159 ,id_160 ,id_161 ,id_162 ,id_163 ,id_164 ,id_165 ,id_166 ,id_167 ,id_168 ,id_169 ,id_170 ,id_171 ,id_172 ,id_173 ,id_174 ,id_175 ,id_176 ,id_177 ,id_178 ,id_179 ,id_180 ,id_181 ,id_182 ,id_183 ,id_184 ,id_185 ,id_186 ,id_187 ,id_188 ,id_189 ,id_190 ,id_191 ,id_192 ,id_193 ,id_194 ,id_195 ,id_196 ,id_197 ,id_198 ,id_199 ,id_200 ,id_201 ,id_202 ,id_203 ,id_204 ,id_205 ,id_206 ,id_207 ,id_208 ,id_209 ,id_210 ,id_211 ,id_212 ,id_213 ,id_214 ,id_215 ,id_216 ,id_217 ,id_218 ,id_219 ,id_220 ,id_221 ,id_222 ,id_223 ,id_224 ,id_225 ,id_226 ,id_227 ,id_228 ,id_229 ,id_230 ,id_231 ,id_232 ,id_233 ,id_234 ,id_235 ,id_236 ,id_237 ,id_238 ,id_239 ,id_240 ,id_1197 ,id_1455 ,id_1459 ,id_1462 ,id_1469 ,id_1480 ,id_1486 ,id_1492 ,id_1496 ,id_2204 ,id_2208 ,id_2211 ,id_2218 ,id_2224 ,id_2230 ,id_2236 ,id_2239 ,id_2247 ,id_2253 ,id_2256 ,id_3698 ,id_3701 ,id_3705 ,id_3711 ,id_3717 ,id_3723 ,id_3729 ,id_3737 ,id_3743 ,id_3749 ,id_4393 ,id_4394 ,id_4400 ,id_4405 ,id_4410 ,id_4415 ,id_4420 ,id_4427 ,id_4432 ,id_4437 ,id_4526 ,id_4528 ,id_2 ,id_3 ,id_450 ,id_448 ,id_444 ,id_442 ,id_440 ,id_438 ,id_496 ,id_494 ,id_492 ,id_490 ,id_488 ,id_486 ,id_484 ,id_482 ,id_480 ,id_560 ,id_542 ,id_558 ,id_556 ,id_554 ,id_552 ,id_550 ,id_548 ,id_546 ,id_544 ,id_540 ,id_538 ,id_536 ,id_534 ,id_532 ,id_530 ,id_528 ,id_526 ,id_524 ,id_279 ,id_436 ,id_478 ,id_522 ,id_402 ,id_404 ,id_406 ,id_408 ,id_410 ,id_432 ,id_446 ,id_284 ,id_286 ,id_289 ,id_292 ,id_341 ,id_281 ,id_453 ,id_278 ,id_373 ,id_246 ,id_258 ,id_264 ,id_270 ,id_388 ,id_391 ,id_394 ,id_397 ,id_376 ,id_379 ,id_382 ,id_385 ,id_412 ,id_414 ,id_416 ,id_249 ,id_295 ,id_324 ,id_252 ,id_276 ,id_310 ,id_313 ,id_316 ,id_319 ,id_327 ,id_330 ,id_333 ,id_336 ,id_418 ,id_273 ,id_298 ,id_301 ,id_304 ,id_307 ,id_344 ,id_422 ,id_469 ,id_419 ,id_471 ,id_359 ,id_362 ,id_365 ,id_368 ,id_347 ,id_350 ,id_353 ,id_356 ,id_321 ,id_338 ,id_370 ,id_399  );

input id_1, id_5, id_9, id_12, id_15, id_18, id_23, id_26, id_29, id_32, id_35, id_38, id_41, id_44, id_47, id_50, id_53, id_54, id_55, id_56, id_57, id_58, id_59, id_60, id_61, id_62, id_63, id_64, id_65, id_66, id_69, id_70, id_73, id_74, id_75, id_76, id_77, id_78, id_79, id_80, id_81, id_82, id_83, id_84, id_85, id_86, id_87, id_88, id_89, id_94, id_97, id_100, id_103, id_106, id_109, id_110, id_111, id_112, id_113, id_114, id_115, id_118, id_121, id_124, id_127, id_130, id_133, id_134, id_135, id_138, id_141, id_144, id_147, id_150, id_151, id_152, id_153, id_154, id_155, id_156, id_157, id_158, id_159, id_160, id_161, id_162, id_163, id_164, id_165, id_166, id_167, id_168, id_169, id_170, id_171, id_172, id_173, id_174, id_175, id_176, id_177, id_178, id_179, id_180, id_181, id_182, id_183, id_184, id_185, id_186, id_187, id_188, id_189, id_190, id_191, id_192, id_193, id_194, id_195, id_196, id_197, id_198, id_199, id_200, id_201, id_202, id_203, id_204, id_205, id_206, id_207, id_208, id_209, id_210, id_211, id_212, id_213, id_214, id_215, id_216, id_217, id_218, id_219, id_220, id_221, id_222, id_223, id_224, id_225, id_226, id_227, id_228, id_229, id_230, id_231, id_232, id_233, id_234, id_235, id_236, id_237, id_238, id_239, id_240, id_1197, id_1455, id_1459, id_1462, id_1469, id_1480, id_1486, id_1492, id_1496, id_2204, id_2208, id_2211, id_2218, id_2224, id_2230, id_2236, id_2239, id_2247, id_2253, id_2256, id_3698, id_3701, id_3705, id_3711, id_3717, id_3723, id_3729, id_3737, id_3743, id_3749, id_4393, id_4394, id_4400, id_4405, id_4410, id_4415, id_4420, id_4427, id_4432, id_4437, id_4526, id_4528;

output id_2, id_3, id_450, id_448, id_444, id_442, id_440, id_438, id_496, id_494, id_492, id_490, id_488, id_486, id_484, id_482, id_480, id_560, id_542, id_558, id_556, id_554, id_552, id_550, id_548, id_546, id_544, id_540, id_538, id_536, id_534, id_532, id_530, id_528, id_526, id_524, id_279, id_436, id_478, id_522, id_402, id_404, id_406, id_408, id_410, id_432, id_446, id_284, id_286, id_289, id_292, id_341, id_281, id_453, id_278, id_373, id_246, id_258, id_264, id_270, id_388, id_391, id_394, id_397, id_376, id_379, id_382, id_385, id_412, id_414, id_416, id_249, id_295, id_324, id_252, id_276, id_310, id_313, id_316, id_319, id_327, id_330, id_333, id_336, id_418, id_273, id_298, id_301, id_304, id_307, id_344, id_422, id_469, id_419, id_471, id_359, id_362, id_365, id_368, id_347, id_350, id_353, id_356, id_321, id_338, id_370, id_399;

buf ( id_2, id_1);
buf ( id_3, id_1);
not ( id_400, id_57);
and ( id_1184, id_134, id_133);
buf ( id_450, id_1459);
buf ( id_448, id_1469);
buf ( id_444, id_1480);
buf ( id_442, id_1486);
buf ( id_440, id_1492);
buf ( id_438, id_1496);
and ( id_1501, id_162, id_172, id_188, id_199);
buf ( id_496, id_2208);
buf ( id_494, id_2218);
buf ( id_492, id_2224);
buf ( id_490, id_2230);
buf ( id_488, id_2236);
buf ( id_486, id_2239);
buf ( id_484, id_2247);
buf ( id_482, id_2253);
buf ( id_480, id_2256);
and ( id_2857, id_150, id_184, id_228, id_240);
buf ( id_560, id_3698);
buf ( id_542, id_3701);
buf ( id_558, id_3705);
buf ( id_556, id_3711);
buf ( id_554, id_3717);
buf ( id_552, id_3723);
buf ( id_550, id_3729);
buf ( id_548, id_3737);
buf ( id_546, id_3743);
buf ( id_544, id_3749);
buf ( id_540, id_4393);
buf ( id_538, id_4400);
buf ( id_536, id_4405);
buf ( id_534, id_4410);
buf ( id_532, id_4415);
buf ( id_530, id_4420);
buf ( id_528, id_4427);
buf ( id_526, id_4432);
buf ( id_524, id_4437);
and ( id_4442, id_183, id_182, id_185, id_186);
and ( id_4514, id_210, id_152, id_218, id_230);
not ( id_279, id_15);
not ( id_401, id_5);
buf ( id_573, id_1);
not ( id_574, id_5);
not ( id_575, id_5);
not ( id_1178, id_2236);
not ( id_1186, id_2253);
not ( id_1192, id_2256);
buf ( id_1198, id_38);
buf ( id_1205, id_15);
nand ( id_1206, id_12, id_9);
nand ( id_1207, id_12, id_9);
buf ( id_1210, id_38);
not ( id_1458, id_1455);
not ( id_1461, id_1459);
buf ( id_436, id_1462);
not ( id_1464, id_1462);
not ( id_1471, id_1469);
buf ( id_1475, id_106);
not ( id_1482, id_1480);
not ( id_1488, id_1486);
not ( id_1495, id_1492);
not ( id_1499, id_1496);
not ( id_1500, id_106);
buf ( id_1503, id_18);
buf ( id_1512, id_18);
and ( id_1518, id_4528, id_1492);
buf ( id_1524, id_18);
not ( id_1535, id_18);
nand ( id_1541, id_4528, id_1496);
not ( id_2207, id_2204);
not ( id_2210, id_2208);
buf ( id_478, id_2211);
not ( id_2213, id_2211);
not ( id_2220, id_2218);
not ( id_2226, id_2224);
not ( id_2232, id_2230);
not ( id_2238, id_2236);
not ( id_2241, id_2239);
not ( id_2249, id_2247);
not ( id_2255, id_2253);
not ( id_2258, id_2256);
buf ( id_2828, id_4526);
not ( id_3700, id_3698);
not ( id_3703, id_3701);
not ( id_3707, id_3705);
not ( id_3713, id_3711);
not ( id_3719, id_3717);
not ( id_3725, id_3723);
not ( id_3731, id_3729);
not ( id_3739, id_3737);
not ( id_3745, id_3743);
not ( id_3751, id_3749);
not ( id_4121, id_4393);
buf ( id_522, id_4394);
not ( id_4396, id_4394);
not ( id_4402, id_4400);
not ( id_4407, id_4405);
not ( id_4412, id_4410);
not ( id_4417, id_4415);
not ( id_4422, id_4420);
not ( id_4429, id_4427);
not ( id_4434, id_4432);
not ( id_4439, id_4437);
buf ( id_4833, id_4526);
nand ( id_402, id_400, id_401);
not ( id_404, id_2857);
not ( id_406, id_4514);
not ( id_408, id_4442);
not ( id_410, id_1501);
and ( id_2876, id_2857, id_4514);
and ( id_2878, id_4442, id_1501);
buf ( id_432, id_573);
buf ( id_446, id_1475);
not ( id_1519, id_1518);
and ( id_2871, id_4528, id_1458);
nand ( id_2883, id_4528, id_2207);
and ( id_280, id_1184, id_575);
nand ( id_284, id_1197, id_574);
not ( id_286, id_1205);
nand ( id_289, id_1197, id_574);
nand ( id_292, id_1184, id_575);
not ( id_341, id_1205);
not ( id_4839, id_4833);
buf ( id_572, id_573);
buf ( id_581, id_1206);
buf ( id_587, id_1512);
buf ( id_601, id_1206);
buf ( id_606, id_1512);
buf ( id_650, id_1206);
buf ( id_657, id_1512);
buf ( id_671, id_1207);
buf ( id_678, id_1503);
and ( id_777, id_1541, id_1198);
and ( id_1115, id_1541, id_1198);
buf ( id_1336, id_1512);
buf ( id_1350, id_1503);
not ( id_1477, id_1475);
not ( id_1507, id_1503);
not ( id_1514, id_1512);
not ( id_1530, id_1524);
buf ( id_2259, id_1535);
not ( id_2833, id_2828);
not ( id_2872, id_2871);
buf ( id_2886, id_1207);
buf ( id_2892, id_1503);
buf ( id_2905, id_1207);
buf ( id_2909, id_1503);
buf ( id_3622, id_1524);
buf ( id_3635, id_1524);
buf ( id_3755, id_1535);
buf ( id_4640, id_1524);
buf ( id_4653, id_1524);
buf ( id_4873, id_1541);
buf ( id_4876, id_1198);
buf ( id_4881, id_1488);
buf ( id_4889, id_1482);
buf ( id_4905, id_1471);
buf ( id_4916, id_1198);
buf ( id_4921, id_1464);
buf ( id_5175, id_1541);
buf ( id_5178, id_1198);
buf ( id_5186, id_1198);
buf ( id_5191, id_1488);
buf ( id_5199, id_1482);
buf ( id_5215, id_1471);
buf ( id_5223, id_1464);
buf ( id_5393, id_1192);
buf ( id_5401, id_1186);
buf ( id_5409, id_2249);
buf ( id_5417, id_1178);
buf ( id_5425, id_2232);
buf ( id_5433, id_2226);
buf ( id_5441, id_2220);
buf ( id_5449, id_2241);
buf ( id_5457, id_2213);
buf ( id_5745, id_1192);
buf ( id_5753, id_1186);
buf ( id_5761, id_2249);
buf ( id_5769, id_2241);
buf ( id_5777, id_1178);
buf ( id_5785, id_2232);
buf ( id_5793, id_2226);
buf ( id_5801, id_2220);
buf ( id_5809, id_2213);
buf ( id_5865, id_3751);
buf ( id_5873, id_3745);
buf ( id_5881, id_3739);
buf ( id_5889, id_3731);
buf ( id_5897, id_3725);
buf ( id_5905, id_3719);
buf ( id_5913, id_3713);
buf ( id_5921, id_3707);
buf ( id_5985, id_3751);
buf ( id_5993, id_3745);
buf ( id_6001, id_3739);
buf ( id_6009, id_3725);
buf ( id_6017, id_3719);
buf ( id_6025, id_3713);
buf ( id_6033, id_3707);
buf ( id_6041, id_3731);
buf ( id_6514, id_1210);
buf ( id_6554, id_1210);
buf ( id_6567, id_4439);
buf ( id_6575, id_4434);
buf ( id_6583, id_4429);
buf ( id_6591, id_4422);
buf ( id_6599, id_4417);
buf ( id_6607, id_4412);
buf ( id_6615, id_4407);
buf ( id_6623, id_4402);
buf ( id_6631, id_4396);
buf ( id_6853, id_4439);
buf ( id_6861, id_4434);
buf ( id_6869, id_4429);
buf ( id_6877, id_4417);
buf ( id_6885, id_4412);
buf ( id_6893, id_4407);
buf ( id_6901, id_4402);
buf ( id_6909, id_4422);
buf ( id_6917, id_4396);
not ( id_281, id_280);
buf ( id_453, id_572);
and ( id_784, id_1519, id_1198);
and ( id_1014, id_1198, id_1519);
and ( id_3221, id_2883, id_1210);
buf ( id_4913, id_1519);
buf ( id_5183, id_1519);
nor ( id_5231, id_1198, id_1519);
buf ( id_6511, id_2883);
and ( id_278, id_163, id_572);
buf ( id_615, id_170);
not ( id_594, id_587);
not ( id_611, id_606);
buf ( id_617, id_169);
buf ( id_619, id_168);
buf ( id_621, id_167);
buf ( id_623, id_166);
buf ( id_625, id_165);
buf ( id_627, id_164);
not ( id_664, id_657);
not ( id_685, id_678);
buf ( id_691, id_177);
buf ( id_693, id_176);
buf ( id_695, id_175);
buf ( id_697, id_174);
buf ( id_699, id_173);
buf ( id_701, id_157);
buf ( id_703, id_156);
buf ( id_705, id_155);
buf ( id_707, id_154);
buf ( id_709, id_153);
not ( id_4879, id_4873);
not ( id_4880, id_4876);
not ( id_4887, id_4881);
not ( id_4895, id_4889);
not ( id_4911, id_4905);
not ( id_4927, id_4921);
not ( id_5181, id_5175);
not ( id_5182, id_5178);
not ( id_5190, id_5186);
not ( id_5197, id_5191);
not ( id_5205, id_5199);
not ( id_5221, id_5215);
not ( id_5229, id_5223);
not ( id_1343, id_1336);
not ( id_1357, id_1350);
and ( id_1364, id_181, id_1336);
and ( id_1366, id_171, id_1336);
and ( id_1368, id_180, id_1336);
and ( id_1370, id_179, id_1336);
and ( id_1372, id_178, id_1336);
and ( id_1374, id_161, id_1350);
and ( id_1376, id_151, id_1350);
and ( id_1378, id_160, id_1350);
and ( id_1380, id_159, id_1350);
and ( id_1382, id_158, id_1350);
not ( id_5399, id_5393);
not ( id_5407, id_5401);
not ( id_5415, id_5409);
not ( id_5423, id_5417);
not ( id_5431, id_5425);
not ( id_5439, id_5433);
not ( id_5447, id_5441);
not ( id_5455, id_5449);
not ( id_5463, id_5457);
not ( id_5751, id_5745);
not ( id_5759, id_5753);
not ( id_5767, id_5761);
not ( id_5775, id_5769);
not ( id_5783, id_5777);
not ( id_5791, id_5785);
not ( id_5799, id_5793);
not ( id_5807, id_5801);
not ( id_5815, id_5809);
buf ( id_2019, id_1514);
buf ( id_2032, id_1507);
buf ( id_2117, id_1514);
buf ( id_2130, id_1507);
not ( id_2266, id_2259);
buf ( id_2272, id_1507);
and ( id_2286, id_44, id_2259);
and ( id_2288, id_41, id_2259);
and ( id_2290, id_29, id_2259);
and ( id_2292, id_26, id_2259);
and ( id_2294, id_23, id_2259);
not ( id_5871, id_5865);
not ( id_5879, id_5873);
not ( id_5887, id_5881);
not ( id_5895, id_5889);
not ( id_5903, id_5897);
not ( id_5911, id_5905);
not ( id_5919, id_5913);
not ( id_5927, id_5921);
not ( id_5991, id_5985);
not ( id_5999, id_5993);
not ( id_6007, id_6001);
not ( id_6015, id_6009);
not ( id_6023, id_6017);
not ( id_6031, id_6025);
not ( id_6039, id_6033);
not ( id_6047, id_6041);
not ( id_2899, id_2892);
not ( id_2914, id_2909);
buf ( id_2919, id_209);
buf ( id_2921, id_216);
buf ( id_2923, id_215);
buf ( id_2925, id_214);
buf ( id_2927, id_213);
buf ( id_2929, id_212);
buf ( id_2931, id_211);
and ( id_3173, id_2872, id_1210);
not ( id_6573, id_6567);
not ( id_6581, id_6575);
not ( id_6589, id_6583);
not ( id_6597, id_6591);
not ( id_6605, id_6599);
not ( id_6613, id_6607);
not ( id_6621, id_6615);
not ( id_6629, id_6623);
not ( id_6637, id_6631);
not ( id_3629, id_3622);
not ( id_3642, id_3635);
and ( id_3649, id_1461, id_3622);
and ( id_3651, id_1464, id_3622);
and ( id_3653, id_1471, id_3622);
and ( id_3655, id_1500, id_3622);
and ( id_3657, id_1482, id_3622);
and ( id_3659, id_1488, id_3635);
and ( id_3661, id_1495, id_3635);
and ( id_3663, id_1499, id_3635);
not ( id_3762, id_3755);
buf ( id_3768, id_1507);
and ( id_3782, id_47, id_3755);
and ( id_3784, id_35, id_3755);
and ( id_3786, id_32, id_3755);
and ( id_3788, id_50, id_3755);
and ( id_3790, id_66, id_3755);
not ( id_6859, id_6853);
not ( id_6867, id_6861);
not ( id_6875, id_6869);
not ( id_6883, id_6877);
not ( id_6891, id_6885);
not ( id_6899, id_6893);
not ( id_6907, id_6901);
not ( id_6915, id_6909);
not ( id_6923, id_6917);
buf ( id_4094, id_1530);
buf ( id_4107, id_1530);
buf ( id_4444, id_1530);
buf ( id_4457, id_1530);
not ( id_4647, id_4640);
not ( id_4660, id_4653);
and ( id_4667, id_2210, id_4640);
and ( id_4669, id_2213, id_4640);
and ( id_4671, id_2220, id_4640);
and ( id_4673, id_2226, id_4640);
and ( id_4675, id_2232, id_4640);
and ( id_4677, id_2238, id_4653);
and ( id_4679, id_2241, id_4653);
and ( id_4681, id_2249, id_4653);
and ( id_4683, id_2255, id_4653);
and ( id_4685, id_2258, id_4653);
buf ( id_4897, id_1477);
buf ( id_5207, id_1477);
buf ( id_6551, id_2872);
nand ( id_763, id_4876, id_4879);
nand ( id_764, id_4873, id_4880);
not ( id_886, id_4913);
nand ( id_1005, id_5178, id_5181);
nand ( id_1006, id_5175, id_5182);
not ( id_5189, id_5183);
nand ( id_1018, id_5183, id_5190);
not ( id_5237, id_5231);
not ( id_3169, id_6511);
buf ( id_5239, id_1014);
or ( id_577, id_594, id_615);
or ( id_618, id_594, id_617);
or ( id_620, id_594, id_619);
or ( id_622, id_594, id_621);
or ( id_624, id_611, id_623);
or ( id_626, id_611, id_625);
or ( id_628, id_611, id_627);
or ( id_692, id_664, id_691);
or ( id_694, id_664, id_693);
or ( id_696, id_664, id_695);
or ( id_698, id_664, id_697);
or ( id_700, id_664, id_699);
or ( id_702, id_685, id_701);
or ( id_704, id_685, id_703);
or ( id_706, id_685, id_705);
or ( id_708, id_685, id_707);
or ( id_710, id_685, id_709);
nand ( id_765, id_763, id_764);
not ( id_4903, id_4897);
not ( id_885, id_4916);
nand ( id_1007, id_1005, id_1006);
nand ( id_1017, id_5186, id_5189);
not ( id_5213, id_5207);
and ( id_1363, id_141, id_1343);
and ( id_1365, id_147, id_1343);
and ( id_1367, id_138, id_1343);
and ( id_1369, id_144, id_1343);
and ( id_1371, id_135, id_1343);
and ( id_1373, id_141, id_1357);
and ( id_1375, id_147, id_1357);
and ( id_1377, id_138, id_1357);
and ( id_1379, id_144, id_1357);
and ( id_1381, id_135, id_1357);
not ( id_2026, id_2019);
not ( id_2039, id_2032);
and ( id_2046, id_103, id_2019);
and ( id_2048, id_130, id_2019);
and ( id_2050, id_127, id_2019);
and ( id_2052, id_124, id_2019);
and ( id_2054, id_100, id_2019);
and ( id_2056, id_103, id_2032);
and ( id_2058, id_130, id_2032);
and ( id_2060, id_127, id_2032);
and ( id_2062, id_124, id_2032);
and ( id_2064, id_100, id_2032);
not ( id_2124, id_2117);
not ( id_2137, id_2130);
and ( id_2144, id_115, id_2117);
and ( id_2146, id_118, id_2117);
and ( id_2148, id_97, id_2117);
and ( id_2150, id_94, id_2117);
and ( id_2152, id_121, id_2117);
and ( id_2154, id_115, id_2130);
and ( id_2156, id_118, id_2130);
and ( id_2158, id_97, id_2130);
and ( id_2160, id_94, id_2130);
and ( id_2162, id_121, id_2130);
not ( id_2279, id_2272);
and ( id_2285, id_208, id_2266);
and ( id_2287, id_198, id_2266);
and ( id_2289, id_207, id_2266);
and ( id_2291, id_206, id_2266);
and ( id_2293, id_205, id_2266);
and ( id_2296, id_44, id_2272);
and ( id_2298, id_41, id_2272);
and ( id_2300, id_29, id_2272);
and ( id_2302, id_26, id_2272);
and ( id_2304, id_23, id_2272);
or ( id_2920, id_2899, id_2919);
or ( id_2922, id_2899, id_2921);
or ( id_2924, id_2899, id_2923);
or ( id_2926, id_2899, id_2925);
or ( id_2928, id_2914, id_2927);
or ( id_2930, id_2914, id_2929);
or ( id_2932, id_2914, id_2931);
not ( id_3168, id_6514);
not ( id_3211, id_6551);
and ( id_3648, id_114, id_3629);
and ( id_3650, id_113, id_3629);
and ( id_3652, id_111, id_3629);
and ( id_3654, id_87, id_3629);
and ( id_3656, id_112, id_3629);
and ( id_3658, id_88, id_3642);
and ( id_3660, id_1455, id_3642);
and ( id_3662, id_2204, id_3642);
buf ( id_3665, id_3703);
buf ( id_3666, id_70);
not ( id_3775, id_3768);
and ( id_3781, id_193, id_3762);
and ( id_3783, id_192, id_3762);
and ( id_3785, id_191, id_3762);
and ( id_3787, id_190, id_3762);
and ( id_3789, id_189, id_3762);
and ( id_3792, id_47, id_3768);
and ( id_3794, id_35, id_3768);
and ( id_3796, id_32, id_3768);
and ( id_3798, id_50, id_3768);
and ( id_3800, id_66, id_3768);
not ( id_4101, id_4094);
not ( id_4114, id_4107);
and ( id_4123, id_58, id_4094);
and ( id_4126, id_77, id_4094);
and ( id_4129, id_78, id_4094);
and ( id_4132, id_59, id_4094);
and ( id_4135, id_81, id_4094);
and ( id_4138, id_80, id_4107);
and ( id_4141, id_79, id_4107);
and ( id_4144, id_60, id_4107);
and ( id_4147, id_61, id_4107);
and ( id_4150, id_62, id_4107);
not ( id_4451, id_4444);
not ( id_4464, id_4457);
and ( id_4471, id_69, id_4444);
and ( id_4473, id_70, id_4444);
and ( id_4475, id_74, id_4444);
and ( id_4477, id_76, id_4444);
and ( id_4479, id_75, id_4444);
and ( id_4481, id_73, id_4457);
and ( id_4483, id_53, id_4457);
and ( id_4485, id_54, id_4457);
and ( id_4487, id_55, id_4457);
and ( id_4489, id_56, id_4457);
and ( id_4666, id_82, id_4647);
and ( id_4668, id_65, id_4647);
and ( id_4670, id_83, id_4647);
and ( id_4672, id_84, id_4647);
and ( id_4674, id_85, id_4647);
and ( id_4676, id_64, id_4660);
and ( id_4678, id_63, id_4660);
and ( id_4680, id_86, id_4660);
and ( id_4682, id_109, id_4660);
and ( id_4684, id_110, id_4660);
buf ( id_579, id_577);
buf ( id_629, id_581);
and ( id_633, id_618, id_581);
and ( id_637, id_620, id_581);
and ( id_641, id_622, id_581);
and ( id_645, id_624, id_601);
and ( id_711, id_692, id_650);
and ( id_715, id_694, id_650);
and ( id_719, id_696, id_650);
and ( id_723, id_698, id_650);
and ( id_727, id_700, id_650);
and ( id_731, id_702, id_671);
and ( id_737, id_704, id_671);
and ( id_745, id_706, id_671);
and ( id_751, id_708, id_671);
and ( id_757, id_710, id_671);
nand ( id_887, id_885, id_886);
nand ( id_1019, id_1017, id_1018);
not ( id_5245, id_5239);
or ( id_1383, id_1365, id_1366);
or ( id_1387, id_1367, id_1368);
or ( id_1391, id_1369, id_1370);
or ( id_1395, id_1371, id_1372);
or ( id_1399, id_1375, id_1376);
or ( id_1406, id_1377, id_1378);
or ( id_1412, id_1379, id_1380);
or ( id_1418, id_1381, id_1382);
or ( id_2305, id_2287, id_2288);
or ( id_2308, id_2289, id_2290);
or ( id_2312, id_2291, id_2292);
or ( id_2316, id_2293, id_2294);
and ( id_2933, id_2920, id_2886);
and ( id_2938, id_2922, id_2886);
and ( id_2942, id_2924, id_2886);
and ( id_2946, id_2926, id_2886);
and ( id_2950, id_2928, id_2905);
nand ( id_3170, id_3168, id_3169);
not ( id_3210, id_6554);
or ( id_3667, id_3650, id_3651);
or ( id_3670, id_3652, id_3653);
or ( id_3673, id_3654, id_3655);
or ( id_3676, id_3656, id_3657);
or ( id_3679, id_3658, id_3659);
or ( id_3682, id_3665, id_3635);
or ( id_3686, id_3666, id_3635);
or ( id_3801, id_3781, id_3782);
or ( id_3804, id_3783, id_3784);
or ( id_3807, id_3785, id_3786);
or ( id_3810, id_3787, id_3788);
or ( id_3813, id_3789, id_3790);
buf ( id_4525, id_2886);
or ( id_4686, id_4668, id_4669);
or ( id_4689, id_4670, id_4671);
or ( id_4692, id_4672, id_4673);
or ( id_4695, id_4674, id_4675);
or ( id_4698, id_4676, id_4677);
or ( id_4701, id_4678, id_4679);
or ( id_4704, id_4680, id_4681);
or ( id_4707, id_4682, id_4683);
or ( id_4710, id_4684, id_4685);
and ( id_5271, id_2932, id_2905);
and ( id_5274, id_2930, id_2905);
and ( id_5305, id_628, id_601);
and ( id_5308, id_626, id_601);
or ( id_5318, id_1373, id_1374);
or ( id_6690, id_3648, id_3649);
or ( id_6711, id_3662, id_3663);
or ( id_6714, id_3660, id_3661);
or ( id_7252, id_2285, id_2286);
or ( id_7296, id_1363, id_1364);
or ( id_7466, id_4666, id_4667);
buf ( id_907, id_784);
buf ( id_913, id_784);
buf ( id_1116, id_1014);
and ( id_2045, id_204, id_2026);
and ( id_2047, id_203, id_2026);
and ( id_2049, id_202, id_2026);
and ( id_2051, id_201, id_2026);
and ( id_2053, id_200, id_2026);
and ( id_2055, id_235, id_2039);
and ( id_2057, id_234, id_2039);
and ( id_2059, id_233, id_2039);
and ( id_2061, id_232, id_2039);
and ( id_2063, id_231, id_2039);
and ( id_2143, id_197, id_2124);
and ( id_2145, id_187, id_2124);
and ( id_2147, id_196, id_2124);
and ( id_2149, id_195, id_2124);
and ( id_2151, id_194, id_2124);
and ( id_2153, id_227, id_2137);
and ( id_2155, id_217, id_2137);
and ( id_2157, id_226, id_2137);
and ( id_2159, id_225, id_2137);
and ( id_2161, id_224, id_2137);
and ( id_2295, id_239, id_2279);
and ( id_2297, id_229, id_2279);
and ( id_2299, id_238, id_2279);
and ( id_2301, id_237, id_2279);
and ( id_2303, id_236, id_2279);
nand ( id_3212, id_3210, id_3211);
and ( id_3791, id_223, id_3775);
and ( id_3793, id_222, id_3775);
and ( id_3795, id_221, id_3775);
and ( id_3797, id_220, id_3775);
and ( id_3799, id_219, id_3775);
and ( id_4122, id_4121, id_4101);
and ( id_4125, id_4396, id_4101);
and ( id_4128, id_4402, id_4101);
and ( id_4131, id_4407, id_4101);
and ( id_4134, id_4412, id_4101);
and ( id_4137, id_4417, id_4114);
and ( id_4140, id_4422, id_4114);
and ( id_4143, id_4429, id_4114);
and ( id_4146, id_4434, id_4114);
and ( id_4149, id_4439, id_4114);
and ( id_4470, id_3700, id_4451);
and ( id_4472, id_3703, id_4451);
and ( id_4474, id_3707, id_4451);
and ( id_4476, id_3713, id_4451);
and ( id_4478, id_3719, id_4451);
and ( id_4480, id_3725, id_4464);
and ( id_4482, id_3731, id_4464);
and ( id_4484, id_3739, id_4464);
and ( id_4486, id_3745, id_4464);
and ( id_4488, id_3751, id_4464);
buf ( id_4962, id_765);
buf ( id_5003, id_765);
buf ( id_5234, id_1007);
buf ( id_5242, id_1007);
not ( id_5250, id_4525);
not ( id_5284, id_579);
and ( id_802, id_1488, id_2950);
and ( id_821, id_1482, id_2946);
and ( id_845, id_1477, id_2942);
and ( id_868, id_1471, id_2938);
and ( id_877, id_1464, id_2933);
and ( id_902, id_887, id_765);
or ( id_908, id_777, id_907);
not ( id_1023, id_1019);
and ( id_1035, id_1488, id_2950);
and ( id_1050, id_1482, id_2946);
and ( id_1068, id_1477, id_2942);
and ( id_1086, id_1471, id_2938);
and ( id_1102, id_1464, id_2933);
and ( id_1108, id_1019, id_1007);
or ( id_1117, id_1115, id_1116);
not ( id_5322, id_5318);
and ( id_1553, id_1192, id_757);
and ( id_1567, id_1186, id_751);
and ( id_1584, id_2249, id_745);
and ( id_1590, id_2241, id_737);
and ( id_1606, id_1178, id_731);
and ( id_1624, id_2232, id_1418);
and ( id_1647, id_2226, id_1412);
and ( id_1669, id_2220, id_1406);
and ( id_1677, id_2213, id_1399);
and ( id_1802, id_1192, id_757);
and ( id_1816, id_1186, id_751);
and ( id_1834, id_2249, id_745);
and ( id_1841, id_737, id_2241);
and ( id_1866, id_1178, id_731);
and ( id_1880, id_2232, id_1418);
and ( id_1897, id_2226, id_1412);
and ( id_1914, id_2220, id_1406);
and ( id_1929, id_2213, id_1399);
or ( id_2065, id_2045, id_2046);
or ( id_2069, id_2047, id_2048);
or ( id_2073, id_2049, id_2050);
or ( id_2077, id_2051, id_2052);
or ( id_2081, id_2053, id_2054);
or ( id_2085, id_2055, id_2056);
or ( id_2091, id_2057, id_2058);
or ( id_2099, id_2059, id_2060);
or ( id_2105, id_2061, id_2062);
or ( id_2111, id_2063, id_2064);
or ( id_2163, id_2145, id_2146);
or ( id_2167, id_2147, id_2148);
or ( id_2171, id_2149, id_2150);
or ( id_2175, id_2151, id_2152);
or ( id_2179, id_2155, id_2156);
or ( id_2186, id_2157, id_2158);
or ( id_2192, id_2159, id_2160);
or ( id_2198, id_2161, id_2162);
or ( id_2320, id_2297, id_2298);
or ( id_2323, id_2299, id_2300);
or ( id_2329, id_2301, id_2302);
or ( id_2335, id_2303, id_2304);
and ( id_2962, id_4710, id_727);
and ( id_2970, id_4707, id_723);
and ( id_2977, id_4704, id_719);
and ( id_2979, id_4701, id_715);
and ( id_2989, id_4698, id_711);
and ( id_2998, id_4695, id_1395);
and ( id_3006, id_4692, id_1391);
and ( id_3013, id_4689, id_1387);
and ( id_3015, id_4686, id_1383);
and ( id_3183, id_3679, id_645);
and ( id_3192, id_3676, id_641);
and ( id_3200, id_3673, id_637);
and ( id_3207, id_3670, id_633);
and ( id_3209, id_3667, id_629);
and ( id_3216, id_3212, id_3170);
buf ( id_3222, id_3173);
not ( id_6694, id_6690);
and ( id_3695, id_1535, id_2305);
or ( id_3816, id_3791, id_3792);
or ( id_3821, id_3793, id_3794);
or ( id_3828, id_3795, id_3796);
or ( id_3833, id_3797, id_3798);
or ( id_3838, id_3799, id_3800);
or ( id_4151, id_4125, id_4126);
or ( id_4154, id_4128, id_4129);
or ( id_4157, id_4131, id_4132);
or ( id_4160, id_4134, id_4135);
or ( id_4163, id_4137, id_4138);
or ( id_4166, id_4140, id_4141);
or ( id_4169, id_4143, id_4144);
or ( id_4172, id_4146, id_4147);
or ( id_4175, id_4149, id_4150);
not ( id_7256, id_7252);
not ( id_7300, id_7296);
or ( id_4490, id_4474, id_4475);
or ( id_4493, id_4476, id_4477);
or ( id_4496, id_4478, id_4479);
or ( id_4499, id_4480, id_4481);
or ( id_4502, id_4482, id_4483);
or ( id_4505, id_4484, id_4485);
or ( id_4508, id_4486, id_4487);
or ( id_4511, id_4488, id_4489);
not ( id_7470, id_7466);
buf ( id_4884, id_2950);
buf ( id_4892, id_2946);
buf ( id_4900, id_2942);
buf ( id_4908, id_2938);
buf ( id_4924, id_2933);
buf ( id_4993, id_887);
nor ( id_5011, id_1464, id_2933);
buf ( id_5194, id_2950);
buf ( id_5202, id_2946);
buf ( id_5210, id_2942);
buf ( id_5218, id_2938);
buf ( id_5226, id_2933);
buf ( id_5247, id_2933);
buf ( id_5255, id_2942);
buf ( id_5258, id_2938);
buf ( id_5263, id_2950);
buf ( id_5266, id_2946);
not ( id_5277, id_5271);
not ( id_5278, id_5274);
buf ( id_5281, id_629);
buf ( id_5289, id_637);
buf ( id_5292, id_633);
buf ( id_5297, id_645);
buf ( id_5300, id_641);
not ( id_5311, id_5305);
not ( id_5312, id_5308);
buf ( id_5315, id_1399);
buf ( id_5323, id_1412);
buf ( id_5326, id_1406);
buf ( id_5331, id_731);
buf ( id_5334, id_1418);
buf ( id_5339, id_745);
buf ( id_5342, id_737);
buf ( id_5349, id_757);
buf ( id_5352, id_751);
buf ( id_5396, id_757);
buf ( id_5404, id_751);
buf ( id_5412, id_745);
buf ( id_5420, id_731);
buf ( id_5428, id_1418);
buf ( id_5436, id_1412);
buf ( id_5444, id_1406);
buf ( id_5452, id_737);
buf ( id_5460, id_1399);
nor ( id_5465, id_2241, id_737);
nor ( id_5581, id_2213, id_1399);
buf ( id_5748, id_757);
buf ( id_5756, id_751);
buf ( id_5764, id_745);
buf ( id_5772, id_737);
buf ( id_5780, id_731);
buf ( id_5788, id_1418);
buf ( id_5796, id_1412);
buf ( id_5804, id_1406);
buf ( id_5812, id_1399);
nor ( id_5849, id_737, id_2241);
buf ( id_5929, id_3682);
buf ( id_6049, id_3682);
buf ( id_6367, id_4710);
buf ( id_6370, id_727);
buf ( id_6375, id_4707);
buf ( id_6378, id_723);
buf ( id_6383, id_4704);
buf ( id_6386, id_719);
buf ( id_6391, id_4698);
buf ( id_6394, id_711);
buf ( id_6399, id_4695);
buf ( id_6402, id_1395);
buf ( id_6407, id_4692);
buf ( id_6410, id_1391);
buf ( id_6415, id_4689);
buf ( id_6418, id_1387);
buf ( id_6423, id_4701);
buf ( id_6426, id_715);
buf ( id_6431, id_4686);
buf ( id_6434, id_1383);
buf ( id_6442, id_3813);
buf ( id_6450, id_3810);
buf ( id_6458, id_3807);
buf ( id_6466, id_3801);
buf ( id_6498, id_3804);
buf ( id_6519, id_3679);
buf ( id_6522, id_645);
buf ( id_6527, id_3676);
buf ( id_6530, id_641);
buf ( id_6535, id_3673);
buf ( id_6538, id_637);
buf ( id_6543, id_3670);
buf ( id_6546, id_633);
buf ( id_6559, id_3667);
buf ( id_6562, id_629);
buf ( id_6687, id_3667);
buf ( id_6695, id_3673);
buf ( id_6698, id_3670);
buf ( id_6703, id_3679);
buf ( id_6706, id_3676);
not ( id_6717, id_6711);
not ( id_6718, id_6714);
or ( id_6724, id_2153, id_2154);
or ( id_6768, id_2295, id_2296);
or ( id_7208, id_2143, id_2144);
buf ( id_7221, id_3801);
buf ( id_7229, id_3807);
buf ( id_7232, id_3804);
buf ( id_7239, id_3813);
buf ( id_7242, id_3810);
buf ( id_7249, id_2305);
buf ( id_7257, id_2312);
buf ( id_7260, id_2308);
buf ( id_7268, id_2316);
buf ( id_7293, id_1383);
buf ( id_7301, id_1391);
buf ( id_7304, id_1387);
buf ( id_7309, id_711);
buf ( id_7312, id_1395);
buf ( id_7317, id_719);
buf ( id_7320, id_715);
buf ( id_7327, id_727);
buf ( id_7330, id_723);
buf ( id_7396, id_2316);
buf ( id_7404, id_2312);
buf ( id_7412, id_2308);
buf ( id_7425, id_3686);
buf ( id_7463, id_4686);
buf ( id_7471, id_4692);
buf ( id_7474, id_4689);
buf ( id_7479, id_4698);
buf ( id_7482, id_4695);
buf ( id_7487, id_4704);
buf ( id_7490, id_4701);
buf ( id_7497, id_4710);
buf ( id_7500, id_4707);
or ( id_7507, id_4472, id_4473);
or ( id_7510, id_4470, id_4471);
or ( id_7554, id_4122, id_4123);
nand ( id_1152, id_5234, id_5237);
not ( id_5238, id_5234);
nand ( id_1156, id_5242, id_5245);
not ( id_5246, id_5242);
not ( id_5288, id_5284);
or ( id_3223, id_3221, id_3222);
buf ( id_4942, id_913);
not ( id_4966, id_4962);
not ( id_5007, id_5003);
nand ( id_5279, id_5274, id_5277);
nand ( id_5280, id_5271, id_5278);
nand ( id_5313, id_5308, id_5311);
nand ( id_5314, id_5305, id_5312);
nand ( id_6719, id_6714, id_6717);
nand ( id_6720, id_6711, id_6718);
nand ( id_790, id_4884, id_4887);
not ( id_4888, id_4884);
nand ( id_803, id_4892, id_4895);
not ( id_4896, id_4892);
nand ( id_825, id_4900, id_4903);
not ( id_4904, id_4900);
nand ( id_851, id_4908, id_4911);
not ( id_4912, id_4908);
nand ( id_893, id_4924, id_4927);
not ( id_4928, id_4924);
not ( id_906, id_902);
nand ( id_1024, id_5194, id_5197);
not ( id_5198, id_5194);
nand ( id_1036, id_5202, id_5205);
not ( id_5206, id_5202);
nand ( id_1053, id_5210, id_5213);
not ( id_5214, id_5210);
nand ( id_1072, id_5218, id_5221);
not ( id_5222, id_5218);
nand ( id_1091, id_5226, id_5229);
not ( id_5230, id_5226);
not ( id_1112, id_1108);
nand ( id_1153, id_5231, id_5238);
nand ( id_1157, id_5239, id_5246);
not ( id_1216, id_5247);
not ( id_5261, id_5255);
not ( id_5262, id_5258);
not ( id_5269, id_5263);
not ( id_5270, id_5266);
not ( id_5287, id_5281);
not ( id_1239, id_5288);
not ( id_5295, id_5289);
not ( id_5296, id_5292);
not ( id_5303, id_5297);
not ( id_5304, id_5300);
not ( id_5321, id_5315);
nand ( id_1262, id_5315, id_5322);
not ( id_5329, id_5323);
not ( id_5330, id_5326);
not ( id_5337, id_5331);
not ( id_5338, id_5334);
nand ( id_1544, id_5396, id_5399);
not ( id_5400, id_5396);
nand ( id_1554, id_5404, id_5407);
not ( id_5408, id_5404);
nand ( id_1571, id_5412, id_5415);
not ( id_5416, id_5412);
nand ( id_1596, id_5420, id_5423);
not ( id_5424, id_5420);
nand ( id_1607, id_5428, id_5431);
not ( id_5432, id_5428);
nand ( id_1628, id_5436, id_5439);
not ( id_5440, id_5436);
nand ( id_1653, id_5444, id_5447);
not ( id_5448, id_5444);
nand ( id_1685, id_5452, id_5455);
not ( id_5456, id_5452);
nand ( id_1693, id_5460, id_5463);
not ( id_5464, id_5460);
nand ( id_1793, id_5748, id_5751);
not ( id_5752, id_5748);
nand ( id_1803, id_5756, id_5759);
not ( id_5760, id_5756);
nand ( id_1820, id_5764, id_5767);
not ( id_5768, id_5764);
nand ( id_1848, id_5772, id_5775);
not ( id_5776, id_5772);
nand ( id_1857, id_5780, id_5783);
not ( id_5784, id_5780);
nand ( id_1867, id_5788, id_5791);
not ( id_5792, id_5788);
nand ( id_1883, id_5796, id_5799);
not ( id_5800, id_5796);
nand ( id_1901, id_5804, id_5807);
not ( id_5808, id_5804);
nand ( id_1919, id_5812, id_5815);
not ( id_5816, id_5812);
not ( id_5855, id_5849);
and ( id_2351, id_3751, id_2111);
and ( id_2366, id_3745, id_2105);
and ( id_2384, id_3739, id_2099);
and ( id_2391, id_2091, id_3731);
and ( id_2417, id_3725, id_2085);
and ( id_2431, id_3719, id_2335);
and ( id_2448, id_3713, id_2329);
and ( id_2465, id_3707, id_2323);
not ( id_5935, id_5929);
and ( id_2597, id_3751, id_2111);
and ( id_2612, id_3745, id_2105);
and ( id_2629, id_3739, id_2099);
and ( id_2635, id_3731, id_2091);
and ( id_2652, id_3725, id_2085);
and ( id_2670, id_3719, id_2335);
and ( id_2693, id_3713, id_2329);
and ( id_2715, id_3707, id_2323);
not ( id_6055, id_6049);
and ( id_3059, id_4175, id_3813);
and ( id_3068, id_4172, id_3810);
and ( id_3076, id_4169, id_3807);
and ( id_3079, id_4166, id_3804);
and ( id_3090, id_4163, id_3801);
and ( id_3099, id_4160, id_2175);
and ( id_3107, id_4157, id_2171);
and ( id_3114, id_4154, id_2167);
and ( id_3116, id_4151, id_2163);
not ( id_3220, id_3216);
and ( id_3292, id_4439, id_3838);
and ( id_3308, id_4434, id_3833);
and ( id_3327, id_4429, id_3828);
and ( id_3335, id_3821, id_4422);
and ( id_3362, id_4417, id_3816);
and ( id_3376, id_4412, id_2198);
and ( id_3393, id_4407, id_2192);
and ( id_3410, id_4402, id_2186);
and ( id_3425, id_4396, id_2179);
not ( id_6693, id_6687);
nand ( id_3503, id_6687, id_6694);
not ( id_6701, id_6695);
not ( id_6702, id_6698);
not ( id_6709, id_6703);
not ( id_6710, id_6706);
not ( id_6728, id_6724);
not ( id_6772, id_6768);
and ( id_3853, id_4439, id_3838);
and ( id_3868, id_4434, id_3833);
and ( id_3885, id_4429, id_3828);
and ( id_3891, id_4422, id_3821);
and ( id_3908, id_4417, id_3816);
and ( id_3926, id_4412, id_2198);
and ( id_3949, id_4407, id_2192);
and ( id_3971, id_4402, id_2186);
and ( id_3979, id_4396, id_2179);
not ( id_7212, id_7208);
not ( id_7227, id_7221);
not ( id_7255, id_7249);
nand ( id_4202, id_7249, id_7256);
not ( id_7263, id_7257);
not ( id_7264, id_7260);
not ( id_7272, id_7268);
not ( id_7299, id_7293);
nand ( id_4225, id_7293, id_7300);
not ( id_7307, id_7301);
not ( id_7308, id_7304);
not ( id_7315, id_7309);
not ( id_7316, id_7312);
and ( id_4297, id_4511, id_2081);
and ( id_4305, id_4508, id_2077);
and ( id_4312, id_4505, id_2073);
and ( id_4314, id_4502, id_2069);
and ( id_4324, id_4499, id_2065);
and ( id_4333, id_4496, id_2316);
and ( id_4341, id_4493, id_2312);
and ( id_4348, id_4490, id_2308);
and ( id_4349, id_3686, id_3695);
and ( id_4389, id_2320, id_1535);
not ( id_7469, id_7463);
nand ( id_4530, id_7463, id_7470);
not ( id_7477, id_7471);
not ( id_7478, id_7474);
not ( id_7485, id_7479);
not ( id_7486, id_7482);
not ( id_7513, id_7507);
not ( id_7514, id_7510);
not ( id_7558, id_7554);
not ( id_5017, id_5011);
buf ( id_5099, id_877);
not ( id_5345, id_5339);
not ( id_5346, id_5342);
not ( id_5355, id_5349);
not ( id_5356, id_5352);
nand ( id_5372, id_5279, id_5280);
nand ( id_5380, id_5313, id_5314);
not ( id_5471, id_5465);
buf ( id_5523, id_1590);
not ( id_5587, id_5581);
buf ( id_5669, id_1677);
buf ( id_5857, id_1841);
buf ( id_5868, id_2111);
buf ( id_5876, id_2105);
buf ( id_5884, id_2099);
buf ( id_5892, id_2091);
buf ( id_5900, id_2085);
buf ( id_5908, id_2335);
buf ( id_5916, id_2329);
buf ( id_5924, id_2323);
nor ( id_5969, id_2091, id_3731);
buf ( id_5988, id_2111);
buf ( id_5996, id_2105);
buf ( id_6004, id_2099);
buf ( id_6012, id_2085);
buf ( id_6020, id_2335);
buf ( id_6028, id_2329);
buf ( id_6036, id_2323);
buf ( id_6044, id_2091);
nor ( id_6057, id_3731, id_2091);
buf ( id_6439, id_4175);
buf ( id_6447, id_4172);
buf ( id_6455, id_4169);
buf ( id_6463, id_4163);
buf ( id_6471, id_4160);
buf ( id_6474, id_2175);
buf ( id_6479, id_4157);
buf ( id_6482, id_2171);
buf ( id_6487, id_4154);
buf ( id_6490, id_2167);
buf ( id_6495, id_4166);
buf ( id_6503, id_4151);
buf ( id_6506, id_2163);
buf ( id_6570, id_3838);
buf ( id_6578, id_3833);
buf ( id_6586, id_3828);
buf ( id_6594, id_3821);
buf ( id_6602, id_3816);
buf ( id_6610, id_2198);
buf ( id_6618, id_2192);
buf ( id_6626, id_2186);
buf ( id_6634, id_2179);
nor ( id_6671, id_3821, id_4422);
buf ( id_6721, id_2179);
buf ( id_6729, id_2192);
buf ( id_6732, id_2186);
buf ( id_6737, id_3816);
buf ( id_6740, id_2198);
buf ( id_6745, id_3828);
buf ( id_6748, id_3821);
buf ( id_6755, id_3838);
buf ( id_6758, id_3833);
buf ( id_6765, id_2320);
buf ( id_6773, id_2329);
buf ( id_6776, id_2323);
buf ( id_6781, id_2085);
buf ( id_6784, id_2335);
buf ( id_6789, id_2099);
buf ( id_6792, id_2091);
buf ( id_6799, id_2111);
buf ( id_6802, id_2105);
nand ( id_6832, id_6719, id_6720);
buf ( id_6856, id_3838);
buf ( id_6864, id_3833);
buf ( id_6872, id_3828);
buf ( id_6880, id_3816);
buf ( id_6888, id_2198);
buf ( id_6896, id_2192);
buf ( id_6904, id_2186);
buf ( id_6912, id_3821);
buf ( id_6920, id_2179);
nor ( id_6925, id_4422, id_3821);
nor ( id_7041, id_4396, id_2179);
buf ( id_7205, id_2163);
buf ( id_7213, id_2171);
buf ( id_7216, id_2167);
buf ( id_7224, id_2175);
not ( id_7235, id_7229);
not ( id_7236, id_7232);
not ( id_7245, id_7239);
not ( id_7246, id_7242);
buf ( id_7265, id_2065);
buf ( id_7273, id_2073);
buf ( id_7276, id_2069);
buf ( id_7283, id_2081);
buf ( id_7286, id_2077);
not ( id_7323, id_7317);
not ( id_7324, id_7320);
not ( id_7333, id_7327);
not ( id_7334, id_7330);
buf ( id_7361, id_4511);
buf ( id_7364, id_2081);
buf ( id_7369, id_4508);
buf ( id_7372, id_2077);
buf ( id_7377, id_4505);
buf ( id_7380, id_2073);
buf ( id_7385, id_4499);
buf ( id_7388, id_2065);
buf ( id_7393, id_4496);
buf ( id_7401, id_4493);
buf ( id_7409, id_4490);
buf ( id_7417, id_4502);
buf ( id_7420, id_2069);
buf ( id_7428, id_3695);
not ( id_7493, id_7487);
not ( id_7494, id_7490);
not ( id_7503, id_7497);
not ( id_7504, id_7500);
buf ( id_7515, id_4493);
buf ( id_7518, id_4490);
buf ( id_7523, id_4499);
buf ( id_7526, id_4496);
buf ( id_7531, id_4505);
buf ( id_7534, id_4502);
buf ( id_7541, id_4511);
buf ( id_7544, id_4508);
buf ( id_7551, id_4151);
buf ( id_7559, id_4157);
buf ( id_7562, id_4154);
buf ( id_7567, id_4163);
buf ( id_7570, id_4160);
buf ( id_7575, id_4169);
buf ( id_7578, id_4166);
buf ( id_7585, id_4175);
buf ( id_7588, id_4172);
not ( id_1176, id_1112);
not ( id_957, id_906);
nand ( id_791, id_4881, id_4888);
nand ( id_804, id_4889, id_4896);
nand ( id_826, id_4897, id_4904);
nand ( id_852, id_4905, id_4912);
nand ( id_894, id_4921, id_4928);
nand ( id_1025, id_5191, id_5198);
nand ( id_1037, id_5199, id_5206);
nand ( id_1054, id_5207, id_5214);
nand ( id_1073, id_5215, id_5222);
nand ( id_1092, id_5223, id_5230);
nand ( id_1154, id_1152, id_1153);
nand ( id_1158, id_1156, id_1157);
not ( id_1215, id_5250);
nand ( id_1224, id_5258, id_5261);
nand ( id_1225, id_5255, id_5262);
nand ( id_1233, id_5266, id_5269);
nand ( id_1234, id_5263, id_5270);
not ( id_1238, id_5287);
nand ( id_1247, id_5292, id_5295);
nand ( id_1248, id_5289, id_5296);
nand ( id_1256, id_5300, id_5303);
nand ( id_1257, id_5297, id_5304);
nand ( id_1261, id_5318, id_5321);
nand ( id_1270, id_5326, id_5329);
nand ( id_1271, id_5323, id_5330);
nand ( id_1279, id_5334, id_5337);
nand ( id_1280, id_5331, id_5338);
nand ( id_1545, id_5393, id_5400);
nand ( id_1555, id_5401, id_5408);
nand ( id_1572, id_5409, id_5416);
nand ( id_1597, id_5417, id_5424);
nand ( id_1608, id_5425, id_5432);
nand ( id_1629, id_5433, id_5440);
nand ( id_1654, id_5441, id_5448);
nand ( id_1686, id_5449, id_5456);
nand ( id_1694, id_5457, id_5464);
nand ( id_1794, id_5745, id_5752);
nand ( id_1804, id_5753, id_5760);
nand ( id_1821, id_5761, id_5768);
nand ( id_1849, id_5769, id_5776);
nand ( id_1858, id_5777, id_5784);
nand ( id_1868, id_5785, id_5792);
nand ( id_1884, id_5793, id_5800);
nand ( id_1902, id_5801, id_5808);
nand ( id_1920, id_5809, id_5816);
not ( id_2954, id_6370);
not ( id_2955, id_6367);
not ( id_2963, id_6378);
not ( id_2964, id_6375);
not ( id_2971, id_6386);
not ( id_2972, id_6383);
not ( id_2980, id_6394);
not ( id_2981, id_6391);
not ( id_2990, id_6402);
not ( id_2991, id_6399);
not ( id_2999, id_6410);
not ( id_3000, id_6407);
not ( id_3007, id_6418);
not ( id_3008, id_6415);
not ( id_3016, id_6426);
not ( id_3017, id_6423);
not ( id_3019, id_6434);
not ( id_3020, id_6431);
not ( id_3174, id_6522);
not ( id_3175, id_6519);
not ( id_3184, id_6530);
not ( id_3185, id_6527);
not ( id_3193, id_6538);
not ( id_3194, id_6535);
not ( id_3201, id_6546);
not ( id_3202, id_6543);
not ( id_3213, id_6562);
not ( id_3214, id_6559);
nand ( id_3502, id_6690, id_6693);
nand ( id_3511, id_6698, id_6701);
nand ( id_3512, id_6695, id_6702);
nand ( id_3520, id_6706, id_6709);
nand ( id_3521, id_6703, id_6710);
nand ( id_4201, id_7252, id_7255);
nand ( id_4210, id_7260, id_7263);
nand ( id_4211, id_7257, id_7264);
nand ( id_4224, id_7296, id_7299);
nand ( id_4233, id_7304, id_7307);
nand ( id_4234, id_7301, id_7308);
nand ( id_4242, id_7312, id_7315);
nand ( id_4243, id_7309, id_7316);
nand ( id_4529, id_7466, id_7469);
nand ( id_4538, id_7474, id_7477);
nand ( id_4539, id_7471, id_7478);
nand ( id_4547, id_7482, id_7485);
nand ( id_4548, id_7479, id_7486);
nand ( id_4552, id_7510, id_7513);
nand ( id_4553, id_7507, id_7514);
not ( id_4946, id_4942);
nand ( id_5347, id_5342, id_5345);
nand ( id_5348, id_5339, id_5346);
nand ( id_5357, id_5352, id_5355);
nand ( id_5358, id_5349, id_5356);
nand ( id_7237, id_7232, id_7235);
nand ( id_7238, id_7229, id_7236);
nand ( id_7247, id_7242, id_7245);
nand ( id_7248, id_7239, id_7246);
nand ( id_7325, id_7320, id_7323);
nand ( id_7326, id_7317, id_7324);
nand ( id_7335, id_7330, id_7333);
nand ( id_7336, id_7327, id_7334);
nand ( id_7495, id_7490, id_7493);
nand ( id_7496, id_7487, id_7494);
nand ( id_7505, id_7500, id_7503);
nand ( id_7506, id_7497, id_7504);
not ( id_3244, id_3220);
nand ( id_792, id_790, id_791);
nand ( id_805, id_803, id_804);
nand ( id_827, id_825, id_826);
nand ( id_853, id_851, id_852);
nand ( id_895, id_893, id_894);
nand ( id_1026, id_1024, id_1025);
nand ( id_1038, id_1036, id_1037);
nand ( id_1055, id_1053, id_1054);
nand ( id_1074, id_1072, id_1073);
nand ( id_1093, id_1091, id_1092);
not ( id_1155, id_1154);
nand ( id_1217, id_1215, id_1216);
nand ( id_1226, id_1224, id_1225);
nand ( id_1235, id_1233, id_1234);
nand ( id_1240, id_1238, id_1239);
nand ( id_1249, id_1247, id_1248);
nand ( id_1258, id_1256, id_1257);
nand ( id_1263, id_1261, id_1262);
nand ( id_1272, id_1270, id_1271);
nand ( id_1281, id_1279, id_1280);
not ( id_5376, id_5372);
not ( id_5384, id_5380);
nand ( id_1546, id_1544, id_1545);
nand ( id_1556, id_1554, id_1555);
nand ( id_1573, id_1571, id_1572);
nand ( id_1598, id_1596, id_1597);
nand ( id_1609, id_1607, id_1608);
nand ( id_1630, id_1628, id_1629);
nand ( id_1655, id_1653, id_1654);
nand ( id_1687, id_1685, id_1686);
nand ( id_1695, id_1693, id_1694);
nand ( id_1795, id_1793, id_1794);
nand ( id_1805, id_1803, id_1804);
nand ( id_1822, id_1820, id_1821);
nand ( id_1850, id_1848, id_1849);
nand ( id_1859, id_1857, id_1858);
nand ( id_1869, id_1867, id_1868);
nand ( id_1885, id_1883, id_1884);
nand ( id_1903, id_1901, id_1902);
nand ( id_1921, id_1919, id_1920);
not ( id_5863, id_5857);
nand ( id_2341, id_5868, id_5871);
not ( id_5872, id_5868);
nand ( id_2352, id_5876, id_5879);
not ( id_5880, id_5876);
nand ( id_2370, id_5884, id_5887);
not ( id_5888, id_5884);
nand ( id_2398, id_5892, id_5895);
not ( id_5896, id_5892);
nand ( id_2407, id_5900, id_5903);
not ( id_5904, id_5900);
nand ( id_2418, id_5908, id_5911);
not ( id_5912, id_5908);
nand ( id_2434, id_5916, id_5919);
not ( id_5920, id_5916);
nand ( id_2452, id_5924, id_5927);
not ( id_5928, id_5924);
and ( id_2481, id_3682, id_4389);
not ( id_5975, id_5969);
nand ( id_2587, id_5988, id_5991);
not ( id_5992, id_5988);
nand ( id_2598, id_5996, id_5999);
not ( id_6000, id_5996);
nand ( id_2616, id_6004, id_6007);
not ( id_6008, id_6004);
nand ( id_2641, id_6012, id_6015);
not ( id_6016, id_6012);
nand ( id_2653, id_6020, id_6023);
not ( id_6024, id_6020);
nand ( id_2674, id_6028, id_6031);
not ( id_6032, id_6028);
nand ( id_2699, id_6036, id_6039);
not ( id_6040, id_6036);
and ( id_2724, id_3682, id_4389);
nand ( id_2732, id_6044, id_6047);
not ( id_6048, id_6044);
nand ( id_2956, id_2954, id_2955);
nand ( id_2965, id_2963, id_2964);
nand ( id_2973, id_2971, id_2972);
nand ( id_2982, id_2980, id_2981);
nand ( id_2992, id_2990, id_2991);
nand ( id_3001, id_2999, id_3000);
nand ( id_3009, id_3007, id_3008);
nand ( id_3018, id_3016, id_3017);
nand ( id_3021, id_3019, id_3020);
not ( id_3051, id_6439);
not ( id_3061, id_6447);
not ( id_3070, id_6455);
not ( id_3081, id_6463);
not ( id_3118, id_6495);
nand ( id_3176, id_3174, id_3175);
nand ( id_3186, id_3184, id_3185);
nand ( id_3195, id_3193, id_3194);
nand ( id_3203, id_3201, id_3202);
nand ( id_3215, id_3213, id_3214);
nand ( id_3281, id_6570, id_6573);
not ( id_6574, id_6570);
nand ( id_3293, id_6578, id_6581);
not ( id_6582, id_6578);
nand ( id_3312, id_6586, id_6589);
not ( id_6590, id_6586);
nand ( id_3342, id_6594, id_6597);
not ( id_6598, id_6594);
nand ( id_3351, id_6602, id_6605);
not ( id_6606, id_6602);
nand ( id_3363, id_6610, id_6613);
not ( id_6614, id_6610);
nand ( id_3379, id_6618, id_6621);
not ( id_6622, id_6618);
nand ( id_3397, id_6626, id_6629);
not ( id_6630, id_6626);
nand ( id_3415, id_6634, id_6637);
not ( id_6638, id_6634);
not ( id_6677, id_6671);
nand ( id_3504, id_3502, id_3503);
nand ( id_3513, id_3511, id_3512);
nand ( id_3522, id_3520, id_3521);
not ( id_6727, id_6721);
nand ( id_3526, id_6721, id_6728);
not ( id_6735, id_6729);
not ( id_6736, id_6732);
not ( id_6743, id_6737);
not ( id_6744, id_6740);
not ( id_6771, id_6765);
nand ( id_3549, id_6765, id_6772);
not ( id_6779, id_6773);
not ( id_6780, id_6776);
not ( id_6787, id_6781);
not ( id_6788, id_6784);
not ( id_6836, id_6832);
nand ( id_3843, id_6856, id_6859);
not ( id_6860, id_6856);
nand ( id_3854, id_6864, id_6867);
not ( id_6868, id_6864);
nand ( id_3872, id_6872, id_6875);
not ( id_6876, id_6872);
nand ( id_3897, id_6880, id_6883);
not ( id_6884, id_6880);
nand ( id_3909, id_6888, id_6891);
not ( id_6892, id_6888);
nand ( id_3930, id_6896, id_6899);
not ( id_6900, id_6896);
nand ( id_3955, id_6904, id_6907);
not ( id_6908, id_6904);
nand ( id_3987, id_6912, id_6915);
not ( id_6916, id_6912);
nand ( id_3995, id_6920, id_6923);
not ( id_6924, id_6920);
not ( id_7211, id_7205);
nand ( id_4179, id_7205, id_7212);
not ( id_7219, id_7213);
not ( id_7220, id_7216);
nand ( id_4196, id_7224, id_7227);
not ( id_7228, id_7224);
nand ( id_4203, id_4201, id_4202);
nand ( id_4212, id_4210, id_4211);
not ( id_7271, id_7265);
nand ( id_4220, id_7265, id_7272);
nand ( id_4226, id_4224, id_4225);
nand ( id_4235, id_4233, id_4234);
nand ( id_4244, id_4242, id_4243);
not ( id_4326, id_7393);
not ( id_4335, id_7401);
not ( id_4343, id_7409);
not ( id_4353, id_7428);
nand ( id_4531, id_4529, id_4530);
nand ( id_4540, id_4538, id_4539);
nand ( id_4549, id_4547, id_4548);
nand ( id_4554, id_4552, id_4553);
not ( id_7521, id_7515);
not ( id_7522, id_7518);
not ( id_7529, id_7523);
not ( id_7530, id_7526);
not ( id_7557, id_7551);
nand ( id_4576, id_7551, id_7558);
not ( id_7565, id_7559);
not ( id_7566, id_7562);
not ( id_7573, id_7567);
not ( id_7574, id_7570);
not ( id_5105, id_5099);
nand ( id_5359, id_5357, id_5358);
nand ( id_5362, id_5347, id_5348);
not ( id_5529, id_5523);
not ( id_5675, id_5669);
buf ( id_5932, id_4389);
buf ( id_5977, id_2391);
buf ( id_6052, id_4389);
not ( id_6063, id_6057);
buf ( id_6115, id_2635);
nor ( id_6173, id_3682, id_4389);
buf ( id_6679, id_3335);
not ( id_6751, id_6745);
not ( id_6752, id_6748);
not ( id_6761, id_6755);
not ( id_6762, id_6758);
not ( id_6795, id_6789);
not ( id_6796, id_6792);
not ( id_6805, id_6799);
not ( id_6806, id_6802);
not ( id_6931, id_6925);
buf ( id_6983, id_3891);
not ( id_7047, id_7041);
buf ( id_7129, id_3979);
not ( id_7279, id_7273);
not ( id_7280, id_7276);
not ( id_7289, id_7283);
not ( id_7290, id_7286);
nand ( id_7337, id_7247, id_7248);
nand ( id_7340, id_7237, id_7238);
nand ( id_7353, id_7335, id_7336);
nand ( id_7356, id_7325, id_7326);
not ( id_7537, id_7531);
not ( id_7538, id_7534);
not ( id_7547, id_7541);
not ( id_7548, id_7544);
not ( id_7581, id_7575);
not ( id_7582, id_7578);
not ( id_7591, id_7585);
not ( id_7592, id_7588);
nand ( id_7595, id_7505, id_7506);
nand ( id_7598, id_7495, id_7496);
nand ( id_2342, id_5865, id_5872);
nand ( id_2353, id_5873, id_5880);
nand ( id_2371, id_5881, id_5888);
nand ( id_2399, id_5889, id_5896);
nand ( id_2408, id_5897, id_5904);
nand ( id_2419, id_5905, id_5912);
nand ( id_2435, id_5913, id_5920);
nand ( id_2453, id_5921, id_5928);
nand ( id_2588, id_5985, id_5992);
nand ( id_2599, id_5993, id_6000);
nand ( id_2617, id_6001, id_6008);
nand ( id_2642, id_6009, id_6016);
nand ( id_2654, id_6017, id_6024);
nand ( id_2675, id_6025, id_6032);
nand ( id_2700, id_6033, id_6040);
nand ( id_2733, id_6041, id_6048);
not ( id_3050, id_6442);
not ( id_3060, id_6450);
not ( id_3069, id_6458);
not ( id_3080, id_6466);
not ( id_3091, id_6474);
not ( id_3092, id_6471);
not ( id_3100, id_6482);
not ( id_3101, id_6479);
not ( id_3108, id_6490);
not ( id_3109, id_6487);
not ( id_3117, id_6498);
not ( id_3120, id_6506);
not ( id_3121, id_6503);
nand ( id_3282, id_6567, id_6574);
nand ( id_3294, id_6575, id_6582);
nand ( id_3313, id_6583, id_6590);
nand ( id_3343, id_6591, id_6598);
nand ( id_3352, id_6599, id_6606);
nand ( id_3364, id_6607, id_6614);
nand ( id_3380, id_6615, id_6622);
nand ( id_3398, id_6623, id_6630);
nand ( id_3416, id_6631, id_6638);
nand ( id_3525, id_6724, id_6727);
nand ( id_3534, id_6732, id_6735);
nand ( id_3535, id_6729, id_6736);
nand ( id_3543, id_6740, id_6743);
nand ( id_3544, id_6737, id_6744);
nand ( id_3548, id_6768, id_6771);
nand ( id_3557, id_6776, id_6779);
nand ( id_3558, id_6773, id_6780);
nand ( id_3566, id_6784, id_6787);
nand ( id_3567, id_6781, id_6788);
nand ( id_3844, id_6853, id_6860);
nand ( id_3855, id_6861, id_6868);
nand ( id_3873, id_6869, id_6876);
nand ( id_3898, id_6877, id_6884);
nand ( id_3910, id_6885, id_6892);
nand ( id_3931, id_6893, id_6900);
nand ( id_3956, id_6901, id_6908);
nand ( id_3988, id_6909, id_6916);
nand ( id_3996, id_6917, id_6924);
nand ( id_4178, id_7208, id_7211);
nand ( id_4187, id_7216, id_7219);
nand ( id_4188, id_7213, id_7220);
nand ( id_4197, id_7221, id_7228);
nand ( id_4219, id_7268, id_7271);
not ( id_4289, id_7364);
not ( id_4290, id_7361);
not ( id_4298, id_7372);
not ( id_4299, id_7369);
not ( id_4306, id_7380);
not ( id_4307, id_7377);
not ( id_4315, id_7388);
not ( id_4316, id_7385);
not ( id_4325, id_7396);
not ( id_4334, id_7404);
not ( id_4342, id_7412);
not ( id_4350, id_7420);
not ( id_4351, id_7417);
not ( id_4354, id_7425);
nand ( id_4561, id_7518, id_7521);
nand ( id_4562, id_7515, id_7522);
nand ( id_4570, id_7526, id_7529);
nand ( id_4571, id_7523, id_7530);
nand ( id_4575, id_7554, id_7557);
nand ( id_4584, id_7562, id_7565);
nand ( id_4585, id_7559, id_7566);
nand ( id_4593, id_7570, id_7573);
nand ( id_4594, id_7567, id_7574);
nand ( id_6753, id_6748, id_6751);
nand ( id_6754, id_6745, id_6752);
nand ( id_6763, id_6758, id_6761);
nand ( id_6764, id_6755, id_6762);
nand ( id_6797, id_6792, id_6795);
nand ( id_6798, id_6789, id_6796);
nand ( id_6807, id_6802, id_6805);
nand ( id_6808, id_6799, id_6806);
nand ( id_7281, id_7276, id_7279);
nand ( id_7282, id_7273, id_7280);
nand ( id_7291, id_7286, id_7289);
nand ( id_7292, id_7283, id_7290);
nand ( id_7539, id_7534, id_7537);
nand ( id_7540, id_7531, id_7538);
nand ( id_7549, id_7544, id_7547);
nand ( id_7550, id_7541, id_7548);
nand ( id_7583, id_7578, id_7581);
nand ( id_7584, id_7575, id_7582);
nand ( id_7593, id_7588, id_7591);
nand ( id_7594, id_7585, id_7592);
not ( id_1856, id_1850);
and ( id_920, id_895, id_853, id_827, id_805, id_792);
and ( id_925, id_792, id_821);
and ( id_926, id_805, id_792, id_845);
and ( id_927, id_827, id_792, id_868, id_805);
and ( id_928, id_853, id_827, id_792, id_877, id_805);
and ( id_937, id_805, id_845);
and ( id_938, id_827, id_868, id_805);
and ( id_939, id_853, id_827, id_877, id_805);
and ( id_940, id_895, id_827, id_805, id_853);
and ( id_941, id_805, id_845);
and ( id_942, id_827, id_868, id_805);
and ( id_943, id_853, id_827, id_877, id_805);
and ( id_944, id_827, id_868);
and ( id_945, id_853, id_827, id_877);
and ( id_946, id_895, id_827, id_853);
and ( id_947, id_827, id_868);
and ( id_948, id_853, id_827, id_877);
and ( id_949, id_853, id_877);
and ( id_956, id_895, id_853);
and ( id_1122, id_1038, id_1093, id_1055, id_1026, id_1074);
and ( id_1125, id_1026, id_1050);
and ( id_1126, id_1038, id_1026, id_1068);
and ( id_1127, id_1055, id_1026, id_1086, id_1038);
and ( id_1128, id_1074, id_1055, id_1026, id_1102, id_1038);
and ( id_1132, id_1038, id_1068);
and ( id_1133, id_1055, id_1086, id_1038);
and ( id_1134, id_1074, id_1055, id_1102, id_1038);
and ( id_1137, id_1086, id_1055);
and ( id_1138, id_1074, id_1055, id_1102);
and ( id_1141, id_1074, id_1102);
not ( id_1221, id_1217);
not ( id_1230, id_1226);
not ( id_1244, id_1240);
not ( id_1253, id_1249);
not ( id_1267, id_1263);
not ( id_1276, id_1272);
buf ( id_1284, id_1235);
buf ( id_1288, id_1235);
buf ( id_1292, id_1258);
buf ( id_1296, id_1258);
buf ( id_1300, id_1281);
buf ( id_1304, id_1281);
and ( id_1702, id_1687, id_1573, id_1556, id_1546);
and ( id_1705, id_1546, id_1567);
and ( id_1706, id_1556, id_1546, id_1584);
and ( id_1707, id_1573, id_1546, id_1590, id_1556);
and ( id_1709, id_1556, id_1584);
and ( id_1710, id_1573, id_1590, id_1556);
and ( id_1711, id_1687, id_1573, id_1556);
and ( id_1712, id_1556, id_1584);
and ( id_1713, id_1573, id_1590, id_1556);
and ( id_1714, id_1573, id_1590);
and ( id_1718, id_1695, id_1655, id_1630, id_1609, id_1598);
and ( id_1722, id_1598, id_1624);
and ( id_1723, id_1609, id_1598, id_1647);
and ( id_1724, id_1630, id_1598, id_1669, id_1609);
and ( id_1725, id_1655, id_1630, id_1598, id_1677, id_1609);
and ( id_1733, id_1609, id_1647);
and ( id_1734, id_1630, id_1669, id_1609);
and ( id_1735, id_1655, id_1630, id_1677, id_1609);
and ( id_1736, id_1695, id_1630, id_1609, id_1655);
and ( id_1737, id_1609, id_1647);
and ( id_1738, id_1630, id_1669, id_1609);
and ( id_1739, id_1655, id_1630, id_1677, id_1609);
and ( id_1740, id_1630, id_1669);
and ( id_1741, id_1655, id_1630, id_1677);
and ( id_1742, id_1695, id_1630, id_1655);
and ( id_1743, id_1630, id_1669);
and ( id_1744, id_1655, id_1630, id_1677);
and ( id_1745, id_1655, id_1677);
and ( id_1749, id_1687, id_1573);
and ( id_1750, id_1695, id_1655);
and ( id_1935, id_1805, id_1850, id_1822, id_1795);
and ( id_1938, id_1795, id_1816);
and ( id_1939, id_1805, id_1795, id_1834);
and ( id_1940, id_1822, id_1795, id_1841, id_1805);
and ( id_1942, id_1805, id_1834);
and ( id_1943, id_1822, id_1841, id_1805);
and ( id_1944, id_1850, id_1822, id_1805);
and ( id_1945, id_1805, id_1834);
and ( id_1946, id_1841, id_1822, id_1805);
and ( id_1947, id_1822, id_1841);
and ( id_1948, id_1850, id_1822);
and ( id_1949, id_1822, id_1841);
and ( id_1950, id_1869, id_1921, id_1885, id_1859, id_1903);
and ( id_1953, id_1859, id_1880);
and ( id_1954, id_1869, id_1859, id_1897);
and ( id_1955, id_1885, id_1859, id_1914, id_1869);
and ( id_1956, id_1903, id_1885, id_1859, id_1929, id_1869);
and ( id_1960, id_1869, id_1897);
and ( id_1961, id_1885, id_1914, id_1869);
and ( id_1962, id_1903, id_1885, id_1929, id_1869);
and ( id_1965, id_1914, id_1885);
and ( id_1966, id_1903, id_1885, id_1929);
and ( id_1969, id_1903, id_1929);
nand ( id_2343, id_2341, id_2342);
nand ( id_2354, id_2352, id_2353);
nand ( id_2372, id_2370, id_2371);
nand ( id_2400, id_2398, id_2399);
nand ( id_2409, id_2407, id_2408);
nand ( id_2420, id_2418, id_2419);
nand ( id_2436, id_2434, id_2435);
nand ( id_2454, id_2452, id_2453);
nand ( id_2470, id_5932, id_5935);
not ( id_5936, id_5932);
not ( id_5983, id_5977);
nand ( id_2589, id_2587, id_2588);
nand ( id_2600, id_2598, id_2599);
nand ( id_2618, id_2616, id_2617);
nand ( id_2643, id_2641, id_2642);
nand ( id_2655, id_2653, id_2654);
nand ( id_2676, id_2674, id_2675);
nand ( id_2701, id_2699, id_2700);
nand ( id_2734, id_2732, id_2733);
nand ( id_2740, id_6052, id_6055);
not ( id_6056, id_6052);
and ( id_3022, id_3018, id_2973, id_2965, id_2956);
and ( id_3025, id_2956, id_2970);
and ( id_3026, id_2965, id_2956, id_2977);
and ( id_3027, id_2973, id_2956, id_2979, id_2965);
and ( id_3029, id_3021, id_3009, id_3001, id_2992, id_2982);
and ( id_3030, id_2982, id_2998);
and ( id_3031, id_2992, id_2982, id_3006);
and ( id_3032, id_3001, id_2982, id_3013, id_2992);
and ( id_3033, id_3009, id_3001, id_2982, id_3015, id_2992);
nand ( id_3052, id_3050, id_3051);
nand ( id_3062, id_3060, id_3061);
nand ( id_3071, id_3069, id_3070);
nand ( id_3082, id_3080, id_3081);
nand ( id_3093, id_3091, id_3092);
nand ( id_3102, id_3100, id_3101);
nand ( id_3110, id_3108, id_3109);
nand ( id_3119, id_3117, id_3118);
nand ( id_3122, id_3120, id_3121);
and ( id_3228, id_3215, id_3203, id_3195, id_3186, id_3176);
and ( id_3231, id_3176, id_3192);
and ( id_3232, id_3186, id_3176, id_3200);
and ( id_3233, id_3195, id_3176, id_3207, id_3186);
and ( id_3234, id_3203, id_3195, id_3176, id_3209, id_3186);
nand ( id_3283, id_3281, id_3282);
nand ( id_3295, id_3293, id_3294);
nand ( id_3314, id_3312, id_3313);
nand ( id_3344, id_3342, id_3343);
nand ( id_3353, id_3351, id_3352);
nand ( id_3365, id_3363, id_3364);
nand ( id_3381, id_3379, id_3380);
nand ( id_3399, id_3397, id_3398);
nand ( id_3417, id_3415, id_3416);
not ( id_6685, id_6679);
not ( id_3508, id_3504);
not ( id_3517, id_3513);
nand ( id_3527, id_3525, id_3526);
nand ( id_3536, id_3534, id_3535);
nand ( id_3545, id_3543, id_3544);
nand ( id_3550, id_3548, id_3549);
nand ( id_3559, id_3557, id_3558);
nand ( id_3568, id_3566, id_3567);
buf ( id_3571, id_3522);
buf ( id_3575, id_3522);
nand ( id_3845, id_3843, id_3844);
nand ( id_3856, id_3854, id_3855);
nand ( id_3874, id_3872, id_3873);
nand ( id_3899, id_3897, id_3898);
nand ( id_3911, id_3909, id_3910);
nand ( id_3932, id_3930, id_3931);
nand ( id_3957, id_3955, id_3956);
nand ( id_3989, id_3987, id_3988);
nand ( id_3997, id_3995, id_3996);
nand ( id_4180, id_4178, id_4179);
nand ( id_4189, id_4187, id_4188);
nand ( id_4198, id_4196, id_4197);
not ( id_4207, id_4203);
not ( id_4216, id_4212);
nand ( id_4221, id_4219, id_4220);
not ( id_4230, id_4226);
not ( id_4239, id_4235);
buf ( id_4263, id_4244);
buf ( id_4267, id_4244);
nand ( id_4291, id_4289, id_4290);
nand ( id_4300, id_4298, id_4299);
nand ( id_4308, id_4306, id_4307);
nand ( id_4317, id_4315, id_4316);
nand ( id_4327, id_4325, id_4326);
nand ( id_4336, id_4334, id_4335);
nand ( id_4344, id_4342, id_4343);
nand ( id_4352, id_4350, id_4351);
nand ( id_4355, id_4353, id_4354);
not ( id_4535, id_4531);
not ( id_4544, id_4540);
not ( id_4558, id_4554);
nand ( id_4563, id_4561, id_4562);
nand ( id_4572, id_4570, id_4571);
nand ( id_4577, id_4575, id_4576);
nand ( id_4586, id_4584, id_4585);
nand ( id_4595, id_4593, id_4594);
buf ( id_4598, id_4549);
buf ( id_4602, id_4549);
buf ( id_4716, id_1921);
buf ( id_4724, id_1859);
buf ( id_4732, id_1869);
buf ( id_4740, id_1885);
buf ( id_4748, id_1903);
buf ( id_4756, id_1093);
buf ( id_4764, id_1026);
buf ( id_4772, id_1038);
buf ( id_4780, id_1055);
buf ( id_4788, id_1074);
buf ( id_5044, id_895);
buf ( id_5054, id_853);
buf ( id_5064, id_792);
buf ( id_5074, id_827);
buf ( id_5084, id_805);
buf ( id_5094, id_805);
buf ( id_5132, id_895);
buf ( id_5142, id_853);
buf ( id_5152, id_792);
buf ( id_5162, id_827);
not ( id_5365, id_5359);
not ( id_5366, id_5362);
buf ( id_5488, id_1687);
buf ( id_5498, id_1573);
buf ( id_5508, id_1546);
buf ( id_5518, id_1556);
buf ( id_5546, id_1687);
buf ( id_5556, id_1573);
buf ( id_5566, id_1546);
buf ( id_5576, id_1556);
buf ( id_5614, id_1695);
buf ( id_5624, id_1655);
buf ( id_5634, id_1598);
buf ( id_5644, id_1630);
buf ( id_5654, id_1609);
buf ( id_5664, id_1609);
buf ( id_5702, id_1695);
buf ( id_5712, id_1655);
buf ( id_5722, id_1598);
buf ( id_5732, id_1630);
buf ( id_5820, id_1795);
buf ( id_5828, id_1795);
buf ( id_5836, id_1805);
buf ( id_5844, id_1805);
buf ( id_5852, id_1822);
buf ( id_5860, id_1822);
not ( id_6121, id_6115);
not ( id_6179, id_6173);
buf ( id_6261, id_2724);
not ( id_7359, id_7353);
not ( id_7360, id_7356);
not ( id_7343, id_7337);
not ( id_7344, id_7340);
nand ( id_6809, id_6763, id_6764);
nand ( id_6812, id_6753, id_6754);
nand ( id_6819, id_6807, id_6808);
nand ( id_6822, id_6797, id_6798);
not ( id_6989, id_6983);
not ( id_7135, id_7129);
nand ( id_7345, id_7291, id_7292);
nand ( id_7348, id_7281, id_7282);
not ( id_7601, id_7595);
not ( id_7602, id_7598);
nand ( id_7603, id_7549, id_7550);
nand ( id_7606, id_7539, id_7540);
nand ( id_7611, id_7593, id_7594);
nand ( id_7614, id_7583, id_7584);
or ( id_929, id_802, id_925, id_926, id_927, id_928);
or ( id_950, id_868, id_949);
or ( id_1129, id_1035, id_1125, id_1126, id_1127, id_1128);
or ( id_1708, id_1553, id_1705, id_1706, id_1707);
or ( id_1715, id_1584, id_1714);
or ( id_1726, id_1606, id_1722, id_1723, id_1724, id_1725);
or ( id_1746, id_1669, id_1745);
or ( id_1941, id_1802, id_1938, id_1939, id_1940);
or ( id_1957, id_1866, id_1953, id_1954, id_1955, id_1956);
nand ( id_2471, id_5929, id_5936);
nand ( id_2741, id_6049, id_6056);
or ( id_3028, id_2962, id_3025, id_3026, id_3027);
or ( id_3034, id_2989, id_3030, id_3031, id_3032, id_3033);
or ( id_3235, id_3183, id_3231, id_3232, id_3233, id_3234);
or ( id_5014, id_845, id_944, id_945, id_946);
or ( id_5034, id_821, id_937, id_938, id_939, id_940);
nor ( id_5102, id_845, id_947, id_948);
nor ( id_5122, id_821, id_941, id_942, id_943);
nand ( id_5367, id_5362, id_5365);
nand ( id_5368, id_5359, id_5366);
or ( id_5478, id_1567, id_1709, id_1710, id_1711);
nor ( id_5536, id_1567, id_1712, id_1713);
or ( id_5584, id_1647, id_1740, id_1741, id_1742);
or ( id_5604, id_1624, id_1733, id_1734, id_1735, id_1736);
nor ( id_5672, id_1647, id_1743, id_1744);
nor ( id_5692, id_1624, id_1737, id_1738, id_1739);
or ( id_5817, id_1816, id_1942, id_1943, id_1944);
nor ( id_5825, id_1816, id_1945, id_1946);
or ( id_5833, id_1834, id_1947, id_1948);
nor ( id_5841, id_1834, id_1949);
nand ( id_6340, id_7356, id_7359);
nand ( id_6341, id_7353, id_7360);
nand ( id_6350, id_7340, id_7343);
nand ( id_6351, id_7337, id_7344);
nand ( id_7436, id_7598, id_7601);
nand ( id_7437, id_7595, id_7602);
not ( id_4720, id_4716);
not ( id_4728, id_4724);
not ( id_4736, id_4732);
not ( id_4744, id_4740);
not ( id_4752, id_4748);
not ( id_4760, id_4756);
not ( id_4768, id_4764);
not ( id_4776, id_4772);
not ( id_4784, id_4780);
not ( id_4792, id_4788);
not ( id_3350, id_3344);
not ( id_2406, id_2400);
not ( id_924, id_920);
not ( id_5088, id_5084);
not ( id_5098, id_5094);
and ( id_997, id_902, id_920);
and ( id_1146, id_1108, id_1122);
not ( id_1287, id_1284);
not ( id_1291, id_1288);
not ( id_1295, id_1292);
not ( id_1299, id_1296);
not ( id_1303, id_1300);
not ( id_1307, id_1304);
and ( id_1309, id_1226, id_1217, id_1284);
and ( id_1312, id_1230, id_1221, id_1288);
and ( id_1315, id_1249, id_1240, id_1292);
and ( id_1318, id_1253, id_1244, id_1296);
and ( id_1321, id_1272, id_1263, id_1300);
and ( id_1324, id_1276, id_1267, id_1304);
not ( id_1721, id_1718);
not ( id_5522, id_5518);
not ( id_5580, id_5576);
not ( id_5658, id_5654);
not ( id_5668, id_5664);
and ( id_1788, id_1702, id_1718);
and ( id_1974, id_1935, id_1950);
not ( id_5824, id_5820);
not ( id_5832, id_5828);
not ( id_5840, id_5836);
not ( id_5848, id_5844);
nand ( id_1999, id_5852, id_5855);
not ( id_5856, id_5852);
nand ( id_2003, id_5860, id_5863);
not ( id_5864, id_5860);
nand ( id_2472, id_2470, id_2471);
and ( id_2487, id_2354, id_2400, id_2372, id_2343);
and ( id_2492, id_2343, id_2366);
and ( id_2493, id_2354, id_2343, id_2384);
and ( id_2494, id_2372, id_2343, id_2391, id_2354);
and ( id_2500, id_2354, id_2384);
and ( id_2501, id_2372, id_2391, id_2354);
and ( id_2502, id_2400, id_2372, id_2354);
and ( id_2503, id_2354, id_2384);
and ( id_2504, id_2391, id_2372, id_2354);
and ( id_2505, id_2372, id_2391);
and ( id_2506, id_2400, id_2372);
and ( id_2507, id_2372, id_2391);
and ( id_2511, id_2409, id_2431);
and ( id_2512, id_2420, id_2409, id_2448);
and ( id_2513, id_2436, id_2409, id_2465, id_2420);
and ( id_2514, id_2454, id_2436, id_2409, id_2481, id_2420);
and ( id_2518, id_2420, id_2448);
and ( id_2519, id_2436, id_2465, id_2420);
and ( id_2520, id_2454, id_2436, id_2481, id_2420);
and ( id_2523, id_2465, id_2436);
and ( id_2524, id_2454, id_2436, id_2481);
and ( id_2527, id_2454, id_2481);
nand ( id_2742, id_2740, id_2741);
and ( id_2749, id_2734, id_2618, id_2600, id_2589);
and ( id_2754, id_2589, id_2612);
and ( id_2755, id_2600, id_2589, id_2629);
and ( id_2756, id_2618, id_2589, id_2635, id_2600);
and ( id_2762, id_2600, id_2629);
and ( id_2763, id_2618, id_2635, id_2600);
and ( id_2764, id_2734, id_2618, id_2600);
and ( id_2765, id_2600, id_2629);
and ( id_2766, id_2618, id_2635, id_2600);
and ( id_2767, id_2618, id_2635);
and ( id_2776, id_2643, id_2670);
and ( id_2777, id_2655, id_2643, id_2693);
and ( id_2778, id_2676, id_2643, id_2715, id_2655);
and ( id_2779, id_2701, id_2676, id_2643, id_2724, id_2655);
and ( id_2788, id_2655, id_2693);
and ( id_2789, id_2676, id_2715, id_2655);
and ( id_2790, id_2701, id_2676, id_2724, id_2655);
and ( id_2792, id_2655, id_2693);
and ( id_2793, id_2676, id_2715, id_2655);
and ( id_2794, id_2701, id_2676, id_2724, id_2655);
and ( id_2795, id_2676, id_2715);
and ( id_2796, id_2701, id_2676, id_2724);
and ( id_2798, id_2676, id_2715);
and ( id_2799, id_2701, id_2676, id_2724);
and ( id_2800, id_2701, id_2724);
and ( id_2804, id_2734, id_2618);
and ( id_3035, id_3022, id_3029);
and ( id_3045, id_3022, id_3034);
and ( id_3123, id_3119, id_3071, id_3062, id_3052);
and ( id_3128, id_3052, id_3068);
and ( id_3129, id_3062, id_3052, id_3076);
and ( id_3130, id_3071, id_3052, id_3079, id_3062);
and ( id_3136, id_3122, id_3110, id_3102, id_3093, id_3082);
and ( id_3139, id_3082, id_3099);
and ( id_3140, id_3093, id_3082, id_3107);
and ( id_3141, id_3102, id_3082, id_3114, id_3093);
and ( id_3142, id_3110, id_3102, id_3082, id_3116, id_3093);
and ( id_3249, id_3216, id_3228);
and ( id_3431, id_3295, id_3344, id_3314, id_3283);
and ( id_3434, id_3283, id_3308);
and ( id_3435, id_3295, id_3283, id_3327);
and ( id_3436, id_3314, id_3283, id_3335, id_3295);
and ( id_3438, id_3295, id_3327);
and ( id_3439, id_3314, id_3335, id_3295);
and ( id_3440, id_3344, id_3314, id_3295);
and ( id_3441, id_3295, id_3327);
and ( id_3442, id_3335, id_3314, id_3295);
and ( id_3443, id_3314, id_3335);
and ( id_3444, id_3344, id_3314);
and ( id_3445, id_3314, id_3335);
and ( id_3446, id_3365, id_3417, id_3381, id_3353, id_3399);
and ( id_3449, id_3353, id_3376);
and ( id_3450, id_3365, id_3353, id_3393);
and ( id_3451, id_3381, id_3353, id_3410, id_3365);
and ( id_3452, id_3399, id_3381, id_3353, id_3425, id_3365);
and ( id_3456, id_3365, id_3393);
and ( id_3457, id_3381, id_3410, id_3365);
and ( id_3458, id_3399, id_3381, id_3425, id_3365);
and ( id_3460, id_3410, id_3381);
and ( id_3461, id_3399, id_3381, id_3425);
and ( id_3463, id_3399, id_3425);
not ( id_3531, id_3527);
not ( id_3540, id_3536);
not ( id_3554, id_3550);
not ( id_3563, id_3559);
not ( id_3574, id_3571);
not ( id_3578, id_3575);
buf ( id_3579, id_3545);
buf ( id_3583, id_3545);
buf ( id_3587, id_3568);
buf ( id_3591, id_3568);
and ( id_3596, id_3513, id_3504, id_3571);
and ( id_3599, id_3517, id_3508, id_3575);
and ( id_4004, id_3989, id_3874, id_3856, id_3845);
and ( id_4007, id_3845, id_3868);
and ( id_4008, id_3856, id_3845, id_3885);
and ( id_4009, id_3874, id_3845, id_3891, id_3856);
and ( id_4011, id_3856, id_3885);
and ( id_4012, id_3874, id_3891, id_3856);
and ( id_4013, id_3989, id_3874, id_3856);
and ( id_4014, id_3856, id_3885);
and ( id_4015, id_3874, id_3891, id_3856);
and ( id_4016, id_3874, id_3891);
and ( id_4020, id_3997, id_3957, id_3932, id_3911, id_3899);
and ( id_4024, id_3899, id_3926);
and ( id_4025, id_3911, id_3899, id_3949);
and ( id_4026, id_3932, id_3899, id_3971, id_3911);
and ( id_4027, id_3957, id_3932, id_3899, id_3979, id_3911);
and ( id_4035, id_3911, id_3949);
and ( id_4036, id_3932, id_3971, id_3911);
and ( id_4037, id_3957, id_3932, id_3979, id_3911);
and ( id_4038, id_3997, id_3932, id_3911, id_3957);
and ( id_4039, id_3911, id_3949);
and ( id_4040, id_3932, id_3971, id_3911);
and ( id_4041, id_3957, id_3932, id_3979, id_3911);
and ( id_4042, id_3932, id_3971);
and ( id_4043, id_3957, id_3932, id_3979);
and ( id_4044, id_3997, id_3932, id_3957);
and ( id_4045, id_3932, id_3971);
and ( id_4046, id_3957, id_3932, id_3979);
and ( id_4047, id_3957, id_3979);
and ( id_4051, id_3989, id_3874);
and ( id_4052, id_3997, id_3957);
not ( id_4184, id_4180);
not ( id_4193, id_4189);
buf ( id_4247, id_4198);
buf ( id_4251, id_4198);
buf ( id_4255, id_4221);
buf ( id_4259, id_4221);
not ( id_4266, id_4263);
not ( id_4270, id_4267);
and ( id_4284, id_4235, id_4226, id_4263);
and ( id_4287, id_4239, id_4230, id_4267);
and ( id_4356, id_4352, id_4308, id_4300, id_4291);
and ( id_4361, id_4291, id_4305);
and ( id_4362, id_4300, id_4291, id_4312);
and ( id_4363, id_4308, id_4291, id_4314, id_4300);
and ( id_4369, id_4355, id_4344, id_4336, id_4327, id_4317);
and ( id_4372, id_4317, id_4333);
and ( id_4373, id_4327, id_4317, id_4341);
and ( id_4374, id_4336, id_4317, id_4348, id_4327);
and ( id_4375, id_4344, id_4336, id_4317, id_4349, id_4327);
not ( id_4567, id_4563);
not ( id_4581, id_4577);
not ( id_4590, id_4586);
not ( id_4601, id_4598);
not ( id_4605, id_4602);
buf ( id_4606, id_4572);
buf ( id_4610, id_4572);
buf ( id_4614, id_4595);
buf ( id_4618, id_4595);
and ( id_4623, id_4540, id_4531, id_4598);
and ( id_4626, id_4544, id_4535, id_4602);
buf ( id_4796, id_3417);
buf ( id_4804, id_3353);
buf ( id_4812, id_3365);
buf ( id_4820, id_3381);
buf ( id_4828, id_3399);
buf ( id_4844, id_2409);
buf ( id_4852, id_2420);
buf ( id_4860, id_2436);
buf ( id_4868, id_2454);
not ( id_4948, id_4946);
not ( id_5048, id_5044);
not ( id_5058, id_5054);
not ( id_5068, id_5064);
not ( id_5078, id_5074);
not ( id_5166, id_5162);
not ( id_5136, id_5132);
not ( id_5146, id_5142);
not ( id_5156, id_5152);
nand ( id_5388, id_5367, id_5368);
not ( id_5492, id_5488);
not ( id_5502, id_5498);
not ( id_5512, id_5508);
not ( id_5550, id_5546);
not ( id_5560, id_5556);
not ( id_5570, id_5566);
not ( id_5618, id_5614);
not ( id_5628, id_5624);
not ( id_5638, id_5634);
not ( id_5648, id_5644);
not ( id_5736, id_5732);
not ( id_5706, id_5702);
not ( id_5716, id_5712);
not ( id_5726, id_5722);
buf ( id_5940, id_2343);
buf ( id_5948, id_2343);
buf ( id_5956, id_2354);
buf ( id_5964, id_2354);
buf ( id_5972, id_2372);
buf ( id_5980, id_2372);
buf ( id_6080, id_2734);
buf ( id_6090, id_2618);
buf ( id_6100, id_2589);
buf ( id_6110, id_2600);
buf ( id_6138, id_2734);
buf ( id_6148, id_2618);
buf ( id_6158, id_2589);
buf ( id_6168, id_2600);
buf ( id_6216, id_2701);
buf ( id_6226, id_2643);
buf ( id_6236, id_2676);
buf ( id_6246, id_2655);
buf ( id_6256, id_2655);
not ( id_6267, id_6261);
buf ( id_6304, id_2701);
buf ( id_6314, id_2643);
buf ( id_6324, id_2676);
nand ( id_6342, id_6340, id_6341);
nand ( id_6352, id_6350, id_6351);
not ( id_7351, id_7345);
not ( id_7352, id_7348);
buf ( id_6642, id_3283);
buf ( id_6650, id_3283);
buf ( id_6658, id_3295);
buf ( id_6666, id_3295);
buf ( id_6674, id_3314);
buf ( id_6682, id_3314);
not ( id_6815, id_6809);
not ( id_6816, id_6812);
not ( id_6825, id_6819);
not ( id_6826, id_6822);
buf ( id_6948, id_3989);
buf ( id_6958, id_3874);
buf ( id_6968, id_3845);
buf ( id_6978, id_3856);
buf ( id_7006, id_3989);
buf ( id_7016, id_3874);
buf ( id_7026, id_3845);
buf ( id_7036, id_3856);
buf ( id_7074, id_3997);
buf ( id_7084, id_3957);
buf ( id_7094, id_3899);
buf ( id_7104, id_3932);
buf ( id_7114, id_3911);
buf ( id_7124, id_3911);
buf ( id_7162, id_3997);
buf ( id_7172, id_3957);
buf ( id_7182, id_3899);
buf ( id_7192, id_3932);
nand ( id_7438, id_7436, id_7437);
not ( id_7617, id_7611);
not ( id_7618, id_7614);
not ( id_7609, id_7603);
not ( id_7610, id_7606);
and ( id_1151, id_1129, id_1108);
and ( id_1002, id_902, id_929);
not ( id_933, id_929);
and ( id_1308, id_1221, id_1226, id_1287);
and ( id_1311, id_1217, id_1230, id_1291);
and ( id_1314, id_1244, id_1249, id_1295);
and ( id_1317, id_1240, id_1253, id_1299);
and ( id_1320, id_1267, id_1272, id_1303);
and ( id_1323, id_1263, id_1276, id_1307);
not ( id_1730, id_1726);
and ( id_1789, id_1702, id_1726);
and ( id_1981, id_1957, id_1935);
not ( id_5823, id_5817);
nand ( id_1986, id_5817, id_5824);
not ( id_5831, id_5825);
nand ( id_1989, id_5825, id_5832);
not ( id_5839, id_5833);
nand ( id_1993, id_5833, id_5840);
not ( id_5847, id_5841);
nand ( id_1996, id_5841, id_5848);
nand ( id_2000, id_5849, id_5856);
nand ( id_2004, id_5857, id_5864);
or ( id_2495, id_2351, id_2492, id_2493, id_2494);
or ( id_2515, id_2417, id_2511, id_2512, id_2513, id_2514);
or ( id_2757, id_2597, id_2754, id_2755, id_2756);
or ( id_2768, id_2629, id_2767);
or ( id_2780, id_2652, id_2776, id_2777, id_2778, id_2779);
or ( id_2801, id_2715, id_2800);
or ( id_3046, id_3028, id_3045);
or ( id_3131, id_3059, id_3128, id_3129, id_3130);
or ( id_3143, id_3090, id_3139, id_3140, id_3141, id_3142);
not ( id_3238, id_3235);
and ( id_3258, id_3216, id_3235);
or ( id_3437, id_3292, id_3434, id_3435, id_3436);
or ( id_3453, id_3362, id_3449, id_3450, id_3451, id_3452);
and ( id_3595, id_3508, id_3513, id_3574);
and ( id_3598, id_3504, id_3517, id_3578);
or ( id_4010, id_3853, id_4007, id_4008, id_4009);
or ( id_4017, id_3885, id_4016);
or ( id_4028, id_3908, id_4024, id_4025, id_4026, id_4027);
or ( id_4048, id_3971, id_4047);
and ( id_4283, id_4230, id_4235, id_4266);
and ( id_4286, id_4226, id_4239, id_4270);
or ( id_4364, id_4297, id_4361, id_4362, id_4363);
or ( id_4376, id_4324, id_4372, id_4373, id_4374, id_4375);
and ( id_4622, id_4535, id_4540, id_4601);
and ( id_4625, id_4531, id_4544, id_4605);
not ( id_5018, id_5014);
nand ( id_5019, id_5014, id_5017);
or ( id_5024, id_950, id_956);
not ( id_5038, id_5034);
not ( id_5106, id_5102);
nand ( id_5107, id_5102, id_5105);
not ( id_5112, id_950);
not ( id_5126, id_5122);
or ( id_5468, id_1715, id_1749);
not ( id_5482, id_5478);
not ( id_5526, id_1715);
not ( id_5540, id_5536);
not ( id_5588, id_5584);
nand ( id_5589, id_5584, id_5587);
or ( id_5594, id_1746, id_1750);
not ( id_5608, id_5604);
not ( id_5676, id_5672);
nand ( id_5677, id_5672, id_5675);
not ( id_5682, id_1746);
not ( id_5696, id_5692);
or ( id_5937, id_2366, id_2500, id_2501, id_2502);
nor ( id_5945, id_2366, id_2503, id_2504);
or ( id_5953, id_2384, id_2505, id_2506);
nor ( id_5961, id_2384, id_2507);
or ( id_6070, id_2612, id_2762, id_2763, id_2764);
nor ( id_6128, id_2612, id_2765, id_2766);
nor ( id_6264, id_2693, id_2798, id_2799);
nor ( id_6284, id_2670, id_2792, id_2793, id_2794);
nand ( id_6360, id_7348, id_7351);
nand ( id_6361, id_7345, id_7352);
or ( id_6639, id_3308, id_3438, id_3439, id_3440);
nor ( id_6647, id_3308, id_3441, id_3442);
or ( id_6655, id_3327, id_3443, id_3444);
nor ( id_6663, id_3327, id_3445);
nand ( id_6817, id_6812, id_6815);
nand ( id_6818, id_6809, id_6816);
nand ( id_6827, id_6822, id_6825);
nand ( id_6828, id_6819, id_6826);
or ( id_6938, id_3868, id_4011, id_4012, id_4013);
nor ( id_6996, id_3868, id_4014, id_4015);
or ( id_7044, id_3949, id_4042, id_4043, id_4044);
or ( id_7064, id_3926, id_4035, id_4036, id_4037, id_4038);
nor ( id_7132, id_3949, id_4045, id_4046);
nor ( id_7152, id_3926, id_4039, id_4040, id_4041);
nand ( id_7446, id_7614, id_7617);
nand ( id_7447, id_7611, id_7618);
nand ( id_7456, id_7606, id_7609);
nand ( id_7457, id_7603, id_7610);
or ( id_241, id_1117, id_1151);
or ( id_265, id_908, id_1002);
nand ( id_2005, id_2003, id_2004);
not ( id_4800, id_4796);
not ( id_4808, id_4804);
not ( id_4816, id_4812);
not ( id_4824, id_4820);
not ( id_4832, id_4828);
not ( id_4848, id_4844);
not ( id_4856, id_4852);
not ( id_4864, id_4860);
not ( id_4872, id_4868);
nor ( id_1310, id_1308, id_1309);
nor ( id_1313, id_1311, id_1312);
nor ( id_1316, id_1314, id_1315);
nor ( id_1319, id_1317, id_1318);
nor ( id_1322, id_1320, id_1321);
nor ( id_1325, id_1323, id_1324);
not ( id_5392, id_5388);
or ( id_1790, id_1708, id_1789);
or ( id_1982, id_1941, id_1981);
nand ( id_1985, id_5820, id_5823);
nand ( id_1988, id_5828, id_5831);
nand ( id_1992, id_5836, id_5839);
nand ( id_1995, id_5844, id_5847);
nand ( id_2001, id_1999, id_2000);
not ( id_2491, id_2487);
and ( id_2508, id_2420, id_2472, id_2436, id_2409, id_2454);
and ( id_2522, id_4526, id_2472, id_2436, id_2454, id_2420);
and ( id_2526, id_4526, id_2472, id_2436, id_2454);
and ( id_2529, id_4526, id_2472, id_2454);
and ( id_2531, id_4526, id_2472);
not ( id_5944, id_5940);
not ( id_5952, id_5948);
not ( id_5960, id_5956);
not ( id_5968, id_5964);
nand ( id_2555, id_5972, id_5975);
not ( id_5976, id_5972);
nand ( id_2559, id_5980, id_5983);
not ( id_5984, id_5980);
not ( id_2753, id_2749);
and ( id_2771, id_2742, id_2701, id_2676, id_2655, id_2643);
and ( id_2791, id_2742, id_2676, id_2655, id_2701);
and ( id_2797, id_2742, id_2676, id_2701);
and ( id_2807, id_2742, id_2701);
not ( id_6114, id_6110);
not ( id_6172, id_6168);
not ( id_6250, id_6246);
not ( id_6260, id_6256);
not ( id_6346, id_6342);
not ( id_6356, id_6352);
not ( id_3127, id_3123);
and ( id_3156, id_3123, id_3136);
or ( id_3259, id_3223, id_3258);
and ( id_3466, id_3431, id_3446);
not ( id_6646, id_6642);
not ( id_6654, id_6650);
not ( id_6662, id_6658);
not ( id_6670, id_6666);
nand ( id_3483, id_6674, id_6677);
not ( id_6678, id_6674);
nand ( id_3487, id_6682, id_6685);
not ( id_6686, id_6682);
not ( id_3582, id_3579);
not ( id_3586, id_3583);
not ( id_3590, id_3587);
not ( id_3594, id_3591);
nor ( id_3597, id_3595, id_3596);
nor ( id_3600, id_3598, id_3599);
and ( id_3602, id_3536, id_3527, id_3579);
and ( id_3605, id_3540, id_3531, id_3583);
and ( id_3608, id_3559, id_3550, id_3587);
and ( id_3611, id_3563, id_3554, id_3591);
not ( id_4023, id_4020);
not ( id_6982, id_6978);
not ( id_7040, id_7036);
not ( id_7118, id_7114);
not ( id_7128, id_7124);
and ( id_4089, id_4004, id_4020);
not ( id_4250, id_4247);
not ( id_4254, id_4251);
not ( id_4258, id_4255);
not ( id_4262, id_4259);
and ( id_4272, id_4189, id_4180, id_4247);
and ( id_4275, id_4193, id_4184, id_4251);
and ( id_4278, id_4212, id_4203, id_4255);
and ( id_4281, id_4216, id_4207, id_4259);
nor ( id_4285, id_4283, id_4284);
nor ( id_4288, id_4286, id_4287);
not ( id_4360, id_4356);
nand ( id_4380, id_4369, id_89);
and ( id_4386, id_4356, id_4369);
not ( id_7442, id_7438);
not ( id_4609, id_4606);
not ( id_4613, id_4610);
not ( id_4617, id_4614);
not ( id_4621, id_4618);
nor ( id_4624, id_4622, id_4623);
nor ( id_4627, id_4625, id_4626);
and ( id_4629, id_4563, id_4554, id_4606);
and ( id_4632, id_4567, id_4558, id_4610);
and ( id_4635, id_4586, id_4577, id_4614);
and ( id_4638, id_4590, id_4581, id_4618);
buf ( id_4836, id_2472);
not ( id_4949, id_4948);
nand ( id_5020, id_5011, id_5018);
nand ( id_5108, id_5099, id_5106);
nand ( id_5590, id_5581, id_5588);
nand ( id_5678, id_5669, id_5676);
not ( id_6084, id_6080);
not ( id_6094, id_6090);
not ( id_6104, id_6100);
not ( id_6142, id_6138);
not ( id_6152, id_6148);
not ( id_6162, id_6158);
buf ( id_6206, id_2742);
not ( id_6220, id_6216);
not ( id_6230, id_6226);
not ( id_6240, id_6236);
not ( id_6328, id_6324);
buf ( id_6294, id_2742);
not ( id_6308, id_6304);
not ( id_6318, id_6314);
nand ( id_6362, id_6360, id_6361);
nand ( id_6840, id_6817, id_6818);
nand ( id_6848, id_6827, id_6828);
not ( id_6952, id_6948);
not ( id_6962, id_6958);
not ( id_6972, id_6968);
not ( id_7010, id_7006);
not ( id_7020, id_7016);
not ( id_7030, id_7026);
not ( id_7078, id_7074);
not ( id_7088, id_7084);
not ( id_7098, id_7094);
not ( id_7108, id_7104);
not ( id_7196, id_7192);
not ( id_7166, id_7162);
not ( id_7176, id_7172);
not ( id_7186, id_7182);
nand ( id_7448, id_7446, id_7447);
nand ( id_7458, id_7456, id_7457);
and ( id_254, id_3046, id_3249);
and ( id_260, id_3046, id_3249);
nand ( id_1987, id_1985, id_1986);
nand ( id_1994, id_1992, id_1993);
not ( id_2002, id_2001);
and ( id_962, id_933, id_924);
and ( id_1751, id_1730, id_1721);
nand ( id_1990, id_1988, id_1989);
nand ( id_1997, id_1995, id_1996);
and ( id_2536, id_2515, id_2487);
not ( id_5943, id_5937);
nand ( id_2542, id_5937, id_5944);
not ( id_5951, id_5945);
nand ( id_2545, id_5945, id_5952);
not ( id_5959, id_5953);
nand ( id_2549, id_5953, id_5960);
not ( id_5967, id_5961);
nand ( id_2552, id_5961, id_5968);
nand ( id_2556, id_5969, id_5976);
nand ( id_2560, id_5977, id_5984);
not ( id_2784, id_2780);
and ( id_2853, id_2749, id_2780);
not ( id_3146, id_3143);
and ( id_3163, id_3123, id_3143);
and ( id_3467, id_3453, id_3431);
not ( id_6645, id_6639);
nand ( id_3470, id_6639, id_6646);
not ( id_6653, id_6647);
nand ( id_3473, id_6647, id_6654);
not ( id_6661, id_6655);
nand ( id_3477, id_6655, id_6662);
not ( id_6669, id_6663);
nand ( id_3480, id_6663, id_6670);
nand ( id_3484, id_6671, id_6678);
nand ( id_3488, id_6679, id_6686);
and ( id_3601, id_3531, id_3536, id_3582);
and ( id_3604, id_3527, id_3540, id_3586);
and ( id_3607, id_3554, id_3559, id_3590);
and ( id_3610, id_3550, id_3563, id_3594);
not ( id_4032, id_4028);
and ( id_4090, id_4004, id_4028);
and ( id_4271, id_4184, id_4189, id_4250);
and ( id_4274, id_4180, id_4193, id_4254);
and ( id_4277, id_4207, id_4212, id_4258);
and ( id_4280, id_4203, id_4216, id_4262);
not ( id_4379, id_4376);
and ( id_4387, id_4356, id_4376);
and ( id_4628, id_4558, id_4563, id_4609);
and ( id_4631, id_4554, id_4567, id_4613);
and ( id_4634, id_4581, id_4586, id_4617);
and ( id_4637, id_4577, id_4590, id_4621);
or ( id_4841, id_2431, id_2518, id_2519, id_2520, id_2522);
or ( id_4849, id_2448, id_2523, id_2524, id_2526);
or ( id_4857, id_2465, id_2527, id_2529);
or ( id_4865, id_2481, id_2531);
nand ( id_5021, id_5019, id_5020);
not ( id_5028, id_5024);
nand ( id_5109, id_5107, id_5108);
not ( id_5116, id_5112);
nand ( id_5369, id_1313, id_1310);
nand ( id_5377, id_1319, id_1316);
nand ( id_5385, id_1325, id_1322);
not ( id_5472, id_5468);
nand ( id_5473, id_5468, id_5471);
not ( id_5530, id_5526);
nand ( id_5531, id_5526, id_5529);
nand ( id_5591, id_5589, id_5590);
not ( id_5598, id_5594);
nand ( id_5679, id_5677, id_5678);
not ( id_5686, id_5682);
or ( id_6060, id_2768, id_2804);
not ( id_6074, id_6070);
not ( id_6118, id_2768);
not ( id_6132, id_6128);
or ( id_6176, id_2693, id_2795, id_2796, id_2797);
or ( id_6186, id_2801, id_2807);
or ( id_6196, id_2670, id_2788, id_2789, id_2790, id_2791);
not ( id_6268, id_6264);
nand ( id_6269, id_6264, id_6267);
not ( id_6274, id_2801);
not ( id_6288, id_6284);
nand ( id_6337, id_4288, id_4285);
nand ( id_6829, id_3600, id_3597);
or ( id_6928, id_4017, id_4051);
not ( id_6942, id_6938);
not ( id_6986, id_4017);
not ( id_7000, id_6996);
not ( id_7048, id_7044);
nand ( id_7049, id_7044, id_7047);
or ( id_7054, id_4048, id_4052);
not ( id_7068, id_7064);
not ( id_7136, id_7132);
nand ( id_7137, id_7132, id_7135);
not ( id_7142, id_4048);
not ( id_7156, id_7152);
nand ( id_7433, id_4627, id_4624);
and ( id_242, id_1982, id_1146);
not ( id_3151, id_3127);
and ( id_257, id_89, id_4386, id_3156, id_3035, id_3249);
and ( id_263, id_89, id_4386, id_3156, id_3035, id_3249);
and ( id_266, id_1790, id_997);
not ( id_1991, id_1990);
not ( id_1998, id_1997);
nand ( id_3489, id_3487, id_3488);
nand ( id_371, id_4836, id_4839);
not ( id_4840, id_4836);
nand ( id_2561, id_2559, id_2560);
and ( id_2532, id_2487, id_2508);
or ( id_2537, id_2495, id_2536);
nand ( id_2541, id_5940, id_5943);
nand ( id_2544, id_5948, id_5951);
nand ( id_2548, id_5956, id_5959);
nand ( id_2551, id_5964, id_5967);
nand ( id_2557, id_2555, id_2556);
and ( id_2563, id_2508, id_4526);
not ( id_2577, id_2491);
not ( id_2775, id_2771);
nand ( id_2806, id_2771, id_4526);
not ( id_2808, id_2753);
and ( id_2852, id_2749, id_2771);
or ( id_2854, id_2757, id_2853);
not ( id_6366, id_6362);
not ( id_4381, id_4360);
or ( id_3164, id_3131, id_3163);
and ( id_3241, id_89, id_4386, id_3156, id_3035);
or ( id_3468, id_3437, id_3467);
nand ( id_3469, id_6642, id_6645);
nand ( id_3472, id_6650, id_6653);
nand ( id_3476, id_6658, id_6661);
nand ( id_3479, id_6666, id_6669);
nand ( id_3485, id_3483, id_3484);
nor ( id_3603, id_3601, id_3602);
nor ( id_3606, id_3604, id_3605);
nor ( id_3609, id_3607, id_3608);
nor ( id_3612, id_3610, id_3611);
not ( id_6844, id_6840);
not ( id_6852, id_6848);
or ( id_4091, id_4010, id_4090);
nor ( id_4273, id_4271, id_4272);
nor ( id_4276, id_4274, id_4275);
nor ( id_4279, id_4277, id_4278);
nor ( id_4282, id_4280, id_4281);
and ( id_4382, id_4379, id_4380);
or ( id_4388, id_4364, id_4387);
not ( id_7452, id_7448);
not ( id_7462, id_7458);
nor ( id_4630, id_4628, id_4629);
nor ( id_4633, id_4631, id_4632);
nor ( id_4636, id_4634, id_4635);
nor ( id_4639, id_4637, id_4638);
not ( id_4958, id_4949);
nand ( id_5474, id_5465, id_5472);
nand ( id_5532, id_5523, id_5530);
not ( id_6210, id_6206);
nand ( id_6270, id_6261, id_6268);
not ( id_6298, id_6294);
nand ( id_7050, id_7041, id_7048);
nand ( id_7138, id_7129, id_7136);
nand ( id_3471, id_3469, id_3470);
nand ( id_3478, id_3476, id_3477);
not ( id_3486, id_3485);
nand ( id_372, id_4833, id_4840);
nand ( id_2543, id_2541, id_2542);
nand ( id_2550, id_2548, id_2549);
not ( id_2558, id_2557);
not ( id_4847, id_4841);
nand ( id_387, id_4841, id_4848);
not ( id_4855, id_4849);
nand ( id_390, id_4849, id_4856);
not ( id_4863, id_4857);
nand ( id_393, id_4857, id_4864);
not ( id_4871, id_4865);
nand ( id_396, id_4865, id_4872);
not ( id_965, id_962);
not ( id_5375, id_5369);
nand ( id_1327, id_5369, id_5376);
not ( id_5383, id_5377);
nand ( id_1330, id_5377, id_5384);
not ( id_5391, id_5385);
nand ( id_1333, id_5385, id_5392);
not ( id_1754, id_1751);
nand ( id_2546, id_2544, id_2545);
nand ( id_2553, id_2551, id_2552);
or ( id_2564, id_2515, id_2563);
and ( id_2809, id_2784, id_2806);
and ( id_2813, id_2784, id_2775);
not ( id_6345, id_6337);
nand ( id_2860, id_6337, id_6346);
nand ( id_3474, id_3472, id_3473);
nand ( id_3481, id_3479, id_3480);
not ( id_6835, id_6829);
nand ( id_3614, id_6829, id_6836);
and ( id_4053, id_4032, id_4023);
not ( id_7441, id_7433);
nand ( id_4516, id_7433, id_7442);
not ( id_4998, id_4993);
not ( id_5027, id_5021);
nand ( id_5030, id_5021, id_5028);
not ( id_5115, id_5109);
nand ( id_5118, id_5109, id_5116);
nand ( id_5475, id_5473, id_5474);
nand ( id_5533, id_5531, id_5532);
not ( id_5597, id_5591);
nand ( id_5600, id_5591, id_5598);
not ( id_5685, id_5679);
nand ( id_5688, id_5679, id_5686);
not ( id_6064, id_6060);
nand ( id_6065, id_6060, id_6063);
not ( id_6122, id_6118);
nand ( id_6123, id_6118, id_6121);
not ( id_6180, id_6176);
nand ( id_6181, id_6176, id_6179);
not ( id_6190, id_6186);
not ( id_6200, id_6196);
nand ( id_6271, id_6269, id_6270);
not ( id_6278, id_6274);
nand ( id_6347, id_4276, id_4273);
nand ( id_6357, id_4282, id_4279);
nand ( id_6837, id_3606, id_3603);
nand ( id_6845, id_3612, id_3609);
not ( id_6932, id_6928);
nand ( id_6933, id_6928, id_6931);
not ( id_6990, id_6986);
nand ( id_6991, id_6986, id_6989);
nand ( id_7051, id_7049, id_7050);
not ( id_7058, id_7054);
nand ( id_7139, id_7137, id_7138);
not ( id_7146, id_7142);
nand ( id_7443, id_4639, id_4636);
nand ( id_7453, id_4633, id_4630);
and ( id_243, id_3468, id_1974, id_1146);
and ( id_244, id_2537, id_3466, id_1974, id_1146);
and ( id_245, id_4526, id_2532, id_3466, id_1974, id_1146);
and ( id_255, id_3164, id_3035, id_3249);
and ( id_256, id_4388, id_3156, id_3035, id_3249);
and ( id_261, id_3164, id_3035, id_3249);
and ( id_262, id_4388, id_3156, id_3035, id_3249);
and ( id_267, id_4091, id_1788, id_997);
and ( id_268, id_2854, id_4089, id_1788, id_997);
and ( id_269, id_4526, id_2852, id_4089, id_1788, id_997);
not ( id_3475, id_3474);
not ( id_3482, id_3481);
nand ( id_373, id_371, id_372);
not ( id_2547, id_2546);
not ( id_2554, id_2553);
nand ( id_386, id_4844, id_4847);
nand ( id_389, id_4852, id_4855);
nand ( id_392, id_4860, id_4863);
nand ( id_395, id_4868, id_4871);
nand ( id_1326, id_5372, id_5375);
nand ( id_1329, id_5380, id_5383);
nand ( id_1332, id_5388, id_5391);
and ( id_1436, id_4091, id_1788);
and ( id_1440, id_2854, id_4089, id_1788);
and ( id_1445, id_4526, id_2852, id_4089, id_1788);
and ( id_1450, id_2854, id_4089);
and ( id_1454, id_4526, id_2852, id_4089);
nand ( id_2859, id_6342, id_6345);
not ( id_4385, id_4382);
buf ( id_3148, id_4364);
and ( id_3239, id_3164, id_3035);
and ( id_3240, id_4388, id_3156, id_3035);
and ( id_3265, id_3468, id_1974);
and ( id_3267, id_2537, id_3466, id_1974);
and ( id_3270, id_4526, id_2532, id_3466, id_1974);
and ( id_3274, id_2537, id_3466);
and ( id_3277, id_4526, id_2532, id_3466);
nand ( id_3613, id_6832, id_6835);
nand ( id_4515, id_7438, id_7441);
not ( id_4959, id_4958);
not ( id_5000, id_4998);
nand ( id_5029, id_5024, id_5027);
nand ( id_5117, id_5112, id_5115);
nand ( id_5599, id_5594, id_5597);
nand ( id_5687, id_5682, id_5685);
nand ( id_6066, id_6057, id_6064);
nand ( id_6124, id_6115, id_6122);
nand ( id_6182, id_6173, id_6180);
nand ( id_6934, id_6925, id_6932);
nand ( id_6992, id_6983, id_6990);
or ( id_246, id_241, id_242, id_243, id_244, id_245);
or ( id_258, id_3259, id_254, id_255, id_256, id_257);
or ( id_264, id_3259, id_260, id_261, id_262, id_263);
or ( id_270, id_265, id_266, id_267, id_268, id_269);
and ( id_375, id_2564, id_2543);
and ( id_378, id_2564, id_2550);
and ( id_381, id_2564, id_2558);
and ( id_384, id_2564, id_2406);
nand ( id_388, id_386, id_387);
nand ( id_391, id_389, id_390);
nand ( id_394, id_392, id_393);
nand ( id_397, id_395, id_396);
nand ( id_1328, id_1326, id_1327);
nand ( id_1331, id_1329, id_1330);
nand ( id_1334, id_1332, id_1333);
or ( id_1447, id_1790, id_1436, id_1440, id_1445);
or ( id_1766, id_4091, id_1450, id_1454);
not ( id_2571, id_2564);
and ( id_2579, id_2577, id_2564);
not ( id_2812, id_2809);
not ( id_2816, id_2813);
buf ( id_2851, id_2757);
nand ( id_2861, id_2859, id_2860);
not ( id_6355, id_6347);
nand ( id_2863, id_6347, id_6356);
not ( id_6365, id_6357);
nand ( id_2866, id_6357, id_6366);
and ( id_3147, id_4381, id_4385);
or ( id_3242, id_3046, id_3239, id_3240, id_3241);
or ( id_3271, id_1982, id_3265, id_3267, id_3270);
or ( id_3279, id_3468, id_3274, id_3277);
nand ( id_3615, id_3613, id_3614);
not ( id_6843, id_6837);
nand ( id_3617, id_6837, id_6844);
not ( id_6851, id_6845);
nand ( id_3620, id_6845, id_6852);
not ( id_4056, id_4053);
nand ( id_4517, id_4515, id_4516);
not ( id_7451, id_7443);
nand ( id_4519, id_7443, id_7452);
not ( id_7461, id_7453);
nand ( id_4522, id_7453, id_7462);
nand ( id_5031, id_5029, id_5030);
nand ( id_5119, id_5117, id_5118);
not ( id_5481, id_5475);
nand ( id_5484, id_5475, id_5482);
not ( id_5539, id_5533);
nand ( id_5542, id_5533, id_5540);
nand ( id_5601, id_5599, id_5600);
nand ( id_5689, id_5687, id_5688);
nand ( id_6067, id_6065, id_6066);
nand ( id_6125, id_6123, id_6124);
nand ( id_6183, id_6181, id_6182);
not ( id_6277, id_6271);
nand ( id_6280, id_6271, id_6278);
nand ( id_6935, id_6933, id_6934);
nand ( id_6993, id_6991, id_6992);
not ( id_7057, id_7051);
nand ( id_7060, id_7051, id_7058);
not ( id_7145, id_7139);
nand ( id_7148, id_7139, id_7146);
nand ( id_4968, id_4959, id_4966);
nand ( id_5009, id_5000, id_5007);
and ( id_2850, id_2808, id_2812);
nand ( id_2862, id_6352, id_6355);
nand ( id_2865, id_6362, id_6365);
or ( id_3149, id_3147, id_3148);
nand ( id_3243, id_3228, id_3242);
nand ( id_3616, id_6840, id_6843);
nand ( id_3619, id_6848, id_6851);
nand ( id_4518, id_7448, id_7451);
nand ( id_4521, id_7458, id_7461);
not ( id_4965, id_4959);
not ( id_5006, id_5000);
nand ( id_5483, id_5478, id_5481);
nand ( id_5541, id_5536, id_5539);
nand ( id_6279, id_6274, id_6277);
nand ( id_7059, id_7054, id_7057);
nand ( id_7147, id_7142, id_7145);
and ( id_374, id_2547, id_2571);
and ( id_377, id_2554, id_2571);
and ( id_380, id_2561, id_2571);
and ( id_383, id_2400, id_2571);
nand ( id_955, id_920, id_1447);
nand ( id_4967, id_4962, id_4965);
nand ( id_5008, id_5003, id_5006);
buf ( id_975, id_1447);
and ( id_1136, id_3271, id_1093, id_1055, id_1074, id_1038);
and ( id_1140, id_3271, id_1093, id_1055, id_1074);
and ( id_1143, id_3271, id_1093, id_1074);
and ( id_1145, id_3271, id_1093);
and ( id_1160, id_1122, id_3271);
not ( id_1771, id_1766);
and ( id_1964, id_3279, id_1921, id_1885, id_1903, id_1869);
and ( id_1968, id_3279, id_1921, id_1885, id_1903);
and ( id_1971, id_3279, id_1921, id_1903);
and ( id_1973, id_3279, id_1921);
and ( id_2007, id_1950, id_3279);
buf ( id_2578, id_2495);
nand ( id_2864, id_2862, id_2863);
nand ( id_2867, id_2865, id_2866);
nand ( id_3150, id_3136, id_3149);
and ( id_3245, id_3238, id_3243);
nand ( id_3618, id_3616, id_3617);
nand ( id_3621, id_3619, id_3620);
or ( id_4067, id_2850, id_2851);
nand ( id_4520, id_4518, id_4519);
nand ( id_4523, id_4521, id_4522);
buf ( id_4713, id_3279);
buf ( id_4753, id_3271);
not ( id_5037, id_5031);
nand ( id_5040, id_5031, id_5038);
not ( id_5125, id_5119);
nand ( id_5128, id_5119, id_5126);
nand ( id_5485, id_5483, id_5484);
nand ( id_5543, id_5541, id_5542);
not ( id_5607, id_5601);
nand ( id_5610, id_5601, id_5608);
not ( id_5695, id_5689);
nand ( id_5698, id_5689, id_5696);
not ( id_6073, id_6067);
nand ( id_6076, id_6067, id_6074);
not ( id_6131, id_6125);
nand ( id_6134, id_6125, id_6132);
not ( id_6189, id_6183);
nand ( id_6192, id_6183, id_6190);
nand ( id_6281, id_6279, id_6280);
not ( id_6941, id_6935);
nand ( id_6944, id_6935, id_6942);
not ( id_6999, id_6993);
nand ( id_7002, id_6993, id_7000);
nand ( id_7061, id_7059, id_7060);
nand ( id_7149, id_7147, id_7148);
or ( id_376, id_374, id_375);
or ( id_379, id_377, id_378);
or ( id_382, id_380, id_381);
or ( id_385, id_383, id_384);
and ( id_958, id_933, id_955);
nand ( id_967, id_4967, id_4968);
nand ( id_971, id_5008, id_5009);
or ( id_1161, id_1129, id_1160);
or ( id_2008, id_1957, id_2007);
or ( id_2580, id_2578, id_2579);
and ( id_2868, id_1331, id_2861, id_2864, id_2867);
and ( id_3152, id_3146, id_3150);
and ( id_4443, id_1328, id_1334, id_3618, id_3621);
and ( id_4524, id_3615, id_4517, id_4520, id_4523);
or ( id_4721, id_1880, id_1960, id_1961, id_1962, id_1964);
or ( id_4729, id_1897, id_1965, id_1966, id_1968);
or ( id_4737, id_1914, id_1969, id_1971);
or ( id_4745, id_1929, id_1973);
or ( id_4761, id_1050, id_1132, id_1133, id_1134, id_1136);
or ( id_4769, id_1068, id_1137, id_1138, id_1140);
or ( id_4777, id_1086, id_1141, id_1143);
or ( id_4785, id_1102, id_1145);
nand ( id_5039, id_5034, id_5037);
nand ( id_5127, id_5122, id_5125);
nand ( id_5609, id_5604, id_5607);
nand ( id_5697, id_5692, id_5695);
nand ( id_6075, id_6070, id_6073);
nand ( id_6133, id_6128, id_6131);
nand ( id_6191, id_6186, id_6189);
nand ( id_6943, id_6938, id_6941);
nand ( id_7001, id_6996, id_6999);
not ( id_3248, id_3245);
buf ( id_248, id_3223);
not ( id_4719, id_4713);
nand ( id_294, id_4713, id_4720);
not ( id_4759, id_4753);
nand ( id_323, id_4753, id_4760);
not ( id_980, id_975);
not ( id_4072, id_4067);
nand ( id_5041, id_5039, id_5040);
nand ( id_5129, id_5127, id_5128);
not ( id_5491, id_5485);
nand ( id_5494, id_5485, id_5492);
not ( id_5549, id_5543);
nand ( id_5552, id_5543, id_5550);
nand ( id_5611, id_5609, id_5610);
nand ( id_5699, id_5697, id_5698);
nand ( id_6077, id_6075, id_6076);
nand ( id_6135, id_6133, id_6134);
nand ( id_6193, id_6191, id_6192);
not ( id_6287, id_6281);
nand ( id_6290, id_6281, id_6288);
nand ( id_6945, id_6943, id_6944);
nand ( id_7003, id_7001, id_7002);
not ( id_7067, id_7061);
nand ( id_7070, id_7061, id_7068);
not ( id_7155, id_7149);
nand ( id_7158, id_7149, id_7156);
and ( id_247, id_3244, id_3248);
not ( id_3155, id_3152);
buf ( id_251, id_3131);
and ( id_272, id_1176, id_1161);
not ( id_961, id_958);
buf ( id_275, id_908);
nand ( id_293, id_4716, id_4719);
and ( id_297, id_2008, id_1987);
and ( id_300, id_2008, id_1994);
and ( id_303, id_2008, id_2002);
and ( id_306, id_2008, id_1856);
not ( id_4727, id_4721);
nand ( id_309, id_4721, id_4728);
not ( id_4735, id_4729);
nand ( id_312, id_4729, id_4736);
not ( id_4743, id_4737);
nand ( id_315, id_4737, id_4744);
not ( id_4751, id_4745);
nand ( id_318, id_4745, id_4752);
nand ( id_322, id_4756, id_4759);
not ( id_4767, id_4761);
nand ( id_326, id_4761, id_4768);
not ( id_4775, id_4769);
nand ( id_329, id_4769, id_4776);
not ( id_4783, id_4777);
nand ( id_332, id_4777, id_4784);
not ( id_4791, id_4785);
nand ( id_335, id_4785, id_4792);
not ( id_412, id_4443);
not ( id_414, id_4524);
not ( id_416, id_2868);
and ( id_2881, id_4443, id_4524, id_2868);
and ( id_993, id_971, id_962);
and ( id_994, id_967, id_965, id_975);
not ( id_1166, id_1161);
and ( id_1171, id_1161, id_1155);
and ( id_1174, id_1161, id_1023);
not ( id_2014, id_2008);
and ( id_3459, id_2580, id_3417, id_3381, id_3399, id_3365);
and ( id_3462, id_2580, id_3417, id_3381, id_3399);
and ( id_3464, id_2580, id_3417, id_3399);
and ( id_3465, id_2580, id_3417);
and ( id_3490, id_3446, id_2580);
buf ( id_4793, id_2580);
nand ( id_5493, id_5488, id_5491);
nand ( id_5551, id_5546, id_5549);
nand ( id_6289, id_6284, id_6287);
nand ( id_7069, id_7064, id_7067);
nand ( id_7157, id_7152, id_7155);
or ( id_249, id_247, id_248);
and ( id_250, id_3151, id_3155);
and ( id_274, id_957, id_961);
nand ( id_295, id_293, id_294);
nand ( id_308, id_4724, id_4727);
nand ( id_311, id_4732, id_4735);
nand ( id_314, id_4740, id_4743);
nand ( id_317, id_4748, id_4751);
nand ( id_324, id_322, id_323);
nand ( id_325, id_4764, id_4767);
nand ( id_328, id_4772, id_4775);
nand ( id_331, id_4780, id_4783);
nand ( id_334, id_4788, id_4791);
and ( id_417, id_2876, id_2878, id_2881);
and ( id_991, id_971, id_933, id_980);
and ( id_992, id_967, id_929);
or ( id_3491, id_3453, id_3490);
or ( id_4801, id_3376, id_3456, id_3457, id_3458, id_3459);
or ( id_4809, id_3393, id_3460, id_3461, id_3462);
or ( id_4817, id_3410, id_3463, id_3464);
or ( id_4825, id_3425, id_3465);
not ( id_5047, id_5041);
nand ( id_5050, id_5041, id_5048);
not ( id_5135, id_5129);
nand ( id_5138, id_5129, id_5136);
nand ( id_5495, id_5493, id_5494);
nand ( id_5553, id_5551, id_5552);
not ( id_5617, id_5611);
nand ( id_5620, id_5611, id_5618);
not ( id_5705, id_5699);
nand ( id_5708, id_5699, id_5706);
not ( id_6083, id_6077);
nand ( id_6086, id_6077, id_6084);
not ( id_6141, id_6135);
nand ( id_6144, id_6135, id_6142);
not ( id_6199, id_6193);
nand ( id_6202, id_6193, id_6200);
nand ( id_6291, id_6289, id_6290);
not ( id_6951, id_6945);
nand ( id_6954, id_6945, id_6952);
not ( id_7009, id_7003);
nand ( id_7012, id_7003, id_7010);
nand ( id_7071, id_7069, id_7070);
nand ( id_7159, id_7157, id_7158);
or ( id_252, id_250, id_251);
buf ( id_271, id_1117);
or ( id_276, id_274, id_275);
and ( id_296, id_1991, id_2014);
and ( id_299, id_1998, id_2014);
and ( id_302, id_2005, id_2014);
and ( id_305, id_1850, id_2014);
nand ( id_310, id_308, id_309);
nand ( id_313, id_311, id_312);
nand ( id_316, id_314, id_315);
nand ( id_319, id_317, id_318);
nand ( id_327, id_325, id_326);
nand ( id_330, id_328, id_329);
nand ( id_333, id_331, id_332);
nand ( id_336, id_334, id_335);
not ( id_4799, id_4793);
nand ( id_343, id_4793, id_4800);
not ( id_418, id_417);
and ( id_1170, id_1158, id_1166);
and ( id_1173, id_1019, id_1166);
nand ( id_5049, id_5044, id_5047);
nand ( id_5137, id_5132, id_5135);
or ( id_5167, id_991, id_992, id_993, id_994);
nand ( id_5619, id_5614, id_5617);
nand ( id_5707, id_5702, id_5705);
nand ( id_6085, id_6080, id_6083);
nand ( id_6143, id_6138, id_6141);
nand ( id_6201, id_6196, id_6199);
nand ( id_6953, id_6948, id_6951);
nand ( id_7011, id_7006, id_7009);
or ( id_273, id_271, id_272);
or ( id_298, id_296, id_297);
or ( id_301, id_299, id_300);
or ( id_304, id_302, id_303);
or ( id_307, id_305, id_306);
nand ( id_342, id_4796, id_4799);
and ( id_346, id_3491, id_3471);
and ( id_349, id_3491, id_3478);
and ( id_352, id_3491, id_3486);
and ( id_355, id_3491, id_3350);
not ( id_4807, id_4801);
nand ( id_358, id_4801, id_4808);
not ( id_4815, id_4809);
nand ( id_361, id_4809, id_4816);
not ( id_4823, id_4817);
nand ( id_364, id_4817, id_4824);
not ( id_4831, id_4825);
nand ( id_367, id_4825, id_4832);
or ( id_1172, id_1170, id_1171);
or ( id_1175, id_1173, id_1174);
not ( id_3497, id_3491);
nand ( id_5051, id_5049, id_5050);
nand ( id_5139, id_5137, id_5138);
not ( id_5501, id_5495);
nand ( id_5504, id_5495, id_5502);
not ( id_5559, id_5553);
nand ( id_5562, id_5553, id_5560);
nand ( id_5621, id_5619, id_5620);
nand ( id_5709, id_5707, id_5708);
nand ( id_6087, id_6085, id_6086);
nand ( id_6145, id_6143, id_6144);
nand ( id_6203, id_6201, id_6202);
not ( id_6297, id_6291);
nand ( id_6300, id_6291, id_6298);
nand ( id_6955, id_6953, id_6954);
nand ( id_7013, id_7011, id_7012);
not ( id_7077, id_7071);
nand ( id_7080, id_7071, id_7078);
not ( id_7165, id_7159);
nand ( id_7168, id_7159, id_7166);
nand ( id_344, id_342, id_343);
nand ( id_357, id_4804, id_4807);
nand ( id_360, id_4812, id_4815);
nand ( id_363, id_4820, id_4823);
nand ( id_366, id_4828, id_4831);
not ( id_5173, id_5167);
buf ( id_422, id_1172);
buf ( id_469, id_1172);
buf ( id_419, id_1175);
buf ( id_471, id_1175);
nand ( id_5503, id_5498, id_5501);
nand ( id_5561, id_5556, id_5559);
nand ( id_6299, id_6294, id_6297);
nand ( id_7079, id_7074, id_7077);
nand ( id_7167, id_7162, id_7165);
and ( id_345, id_3475, id_3497);
and ( id_348, id_3482, id_3497);
and ( id_351, id_3489, id_3497);
and ( id_354, id_3344, id_3497);
nand ( id_359, id_357, id_358);
nand ( id_362, id_360, id_361);
nand ( id_365, id_363, id_364);
nand ( id_368, id_366, id_367);
not ( id_5057, id_5051);
nand ( id_5060, id_5051, id_5058);
not ( id_5145, id_5139);
nand ( id_5148, id_5139, id_5146);
nand ( id_5505, id_5503, id_5504);
nand ( id_5563, id_5561, id_5562);
not ( id_5627, id_5621);
nand ( id_5630, id_5621, id_5628);
not ( id_5715, id_5709);
nand ( id_5718, id_5709, id_5716);
not ( id_6093, id_6087);
nand ( id_6096, id_6087, id_6094);
not ( id_6151, id_6145);
nand ( id_6154, id_6145, id_6152);
not ( id_6209, id_6203);
nand ( id_6212, id_6203, id_6210);
nand ( id_6301, id_6299, id_6300);
not ( id_6961, id_6955);
nand ( id_6964, id_6955, id_6962);
not ( id_7019, id_7013);
nand ( id_7022, id_7013, id_7020);
nand ( id_7081, id_7079, id_7080);
nand ( id_7169, id_7167, id_7168);
or ( id_347, id_345, id_346);
or ( id_350, id_348, id_349);
or ( id_353, id_351, id_352);
or ( id_356, id_354, id_355);
nand ( id_5059, id_5054, id_5057);
nand ( id_5147, id_5142, id_5145);
nand ( id_5629, id_5624, id_5627);
nand ( id_5717, id_5712, id_5715);
nand ( id_6095, id_6090, id_6093);
nand ( id_6153, id_6148, id_6151);
nand ( id_6211, id_6206, id_6209);
nand ( id_6963, id_6958, id_6961);
nand ( id_7021, id_7016, id_7019);
nand ( id_5061, id_5059, id_5060);
nand ( id_5149, id_5147, id_5148);
not ( id_5511, id_5505);
nand ( id_5514, id_5505, id_5512);
not ( id_5569, id_5563);
nand ( id_5572, id_5563, id_5570);
nand ( id_5631, id_5629, id_5630);
nand ( id_5719, id_5717, id_5718);
nand ( id_6097, id_6095, id_6096);
nand ( id_6155, id_6153, id_6154);
nand ( id_6213, id_6211, id_6212);
not ( id_6307, id_6301);
nand ( id_6310, id_6301, id_6308);
nand ( id_6965, id_6963, id_6964);
nand ( id_7023, id_7021, id_7022);
not ( id_7087, id_7081);
nand ( id_7090, id_7081, id_7088);
not ( id_7175, id_7169);
nand ( id_7178, id_7169, id_7176);
nand ( id_5513, id_5508, id_5511);
nand ( id_5571, id_5566, id_5569);
nand ( id_6309, id_6304, id_6307);
nand ( id_7089, id_7084, id_7087);
nand ( id_7177, id_7172, id_7175);
not ( id_5067, id_5061);
nand ( id_5070, id_5061, id_5068);
not ( id_5155, id_5149);
nand ( id_5158, id_5149, id_5156);
nand ( id_5515, id_5513, id_5514);
nand ( id_5573, id_5571, id_5572);
not ( id_5637, id_5631);
nand ( id_5640, id_5631, id_5638);
not ( id_5725, id_5719);
nand ( id_5728, id_5719, id_5726);
not ( id_6103, id_6097);
nand ( id_6106, id_6097, id_6104);
not ( id_6161, id_6155);
nand ( id_6164, id_6155, id_6162);
not ( id_6219, id_6213);
nand ( id_6222, id_6213, id_6220);
nand ( id_6311, id_6309, id_6310);
not ( id_6971, id_6965);
nand ( id_6974, id_6965, id_6972);
not ( id_7029, id_7023);
nand ( id_7032, id_7023, id_7030);
nand ( id_7091, id_7089, id_7090);
nand ( id_7179, id_7177, id_7178);
nand ( id_5069, id_5064, id_5067);
nand ( id_5157, id_5152, id_5155);
nand ( id_5639, id_5634, id_5637);
nand ( id_5727, id_5722, id_5725);
nand ( id_6105, id_6100, id_6103);
nand ( id_6163, id_6158, id_6161);
nand ( id_6221, id_6216, id_6219);
nand ( id_6973, id_6968, id_6971);
nand ( id_7031, id_7026, id_7029);
not ( id_5521, id_5515);
nand ( id_1756, id_5515, id_5522);
not ( id_5579, id_5573);
nand ( id_1761, id_5573, id_5580);
nand ( id_5071, id_5069, id_5070);
nand ( id_5159, id_5157, id_5158);
nand ( id_5641, id_5639, id_5640);
nand ( id_5729, id_5727, id_5728);
nand ( id_6107, id_6105, id_6106);
nand ( id_6165, id_6163, id_6164);
nand ( id_6223, id_6221, id_6222);
not ( id_6317, id_6311);
nand ( id_6320, id_6311, id_6318);
nand ( id_6975, id_6973, id_6974);
nand ( id_7033, id_7031, id_7032);
not ( id_7097, id_7091);
nand ( id_7100, id_7091, id_7098);
not ( id_7185, id_7179);
nand ( id_7188, id_7179, id_7186);
nand ( id_1755, id_5518, id_5521);
nand ( id_1760, id_5576, id_5579);
nand ( id_6319, id_6314, id_6317);
nand ( id_7099, id_7094, id_7097);
nand ( id_7187, id_7182, id_7185);
nand ( id_1757, id_1755, id_1756);
nand ( id_1762, id_1760, id_1761);
not ( id_6113, id_6107);
nand ( id_2818, id_6107, id_6114);
not ( id_6171, id_6165);
nand ( id_2823, id_6165, id_6172);
not ( id_6981, id_6975);
nand ( id_4058, id_6975, id_6982);
not ( id_7039, id_7033);
nand ( id_4063, id_7033, id_7040);
not ( id_5077, id_5071);
nand ( id_5080, id_5071, id_5078);
not ( id_5165, id_5159);
nand ( id_5090, id_5159, id_5166);
not ( id_5647, id_5641);
nand ( id_5650, id_5641, id_5648);
not ( id_5735, id_5729);
nand ( id_5660, id_5729, id_5736);
not ( id_6229, id_6223);
nand ( id_6232, id_6223, id_6230);
nand ( id_6321, id_6319, id_6320);
nand ( id_7101, id_7099, id_7100);
nand ( id_7189, id_7187, id_7188);
nand ( id_2817, id_6110, id_6113);
nand ( id_2822, id_6168, id_6171);
nand ( id_4057, id_6978, id_6981);
nand ( id_4062, id_7036, id_7039);
nand ( id_5079, id_5074, id_5077);
nand ( id_5089, id_5162, id_5165);
nand ( id_5649, id_5644, id_5647);
nand ( id_5659, id_5732, id_5735);
nand ( id_6231, id_6226, id_6229);
and ( id_1782, id_1762, id_1730, id_1771);
and ( id_1783, id_1757, id_1726);
and ( id_1784, id_1762, id_1751);
and ( id_1785, id_1757, id_1754, id_1766);
nand ( id_2819, id_2817, id_2818);
nand ( id_2824, id_2822, id_2823);
nand ( id_4059, id_4057, id_4058);
nand ( id_4064, id_4062, id_4063);
nand ( id_5081, id_5079, id_5080);
nand ( id_5091, id_5089, id_5090);
nand ( id_5651, id_5649, id_5650);
nand ( id_5661, id_5659, id_5660);
nand ( id_6233, id_6231, id_6232);
not ( id_6327, id_6321);
nand ( id_6252, id_6321, id_6328);
not ( id_7107, id_7101);
nand ( id_7110, id_7101, id_7108);
not ( id_7195, id_7189);
nand ( id_7120, id_7189, id_7196);
or ( id_5737, id_1782, id_1783, id_1784, id_1785);
nand ( id_6251, id_6324, id_6327);
nand ( id_7109, id_7104, id_7107);
nand ( id_7119, id_7192, id_7195);
not ( id_5087, id_5081);
nand ( id_985, id_5081, id_5088);
not ( id_5097, id_5091);
nand ( id_988, id_5091, id_5098);
not ( id_5657, id_5651);
nand ( id_1776, id_5651, id_5658);
not ( id_5667, id_5661);
nand ( id_1779, id_5661, id_5668);
and ( id_2844, id_2824, id_2784, id_2833);
and ( id_2845, id_2819, id_2780);
and ( id_2846, id_2824, id_2813);
and ( id_2847, id_2819, id_2816, id_2828);
and ( id_4083, id_4064, id_4032, id_4072);
and ( id_4084, id_4059, id_4028);
and ( id_4085, id_4064, id_4053);
and ( id_4086, id_4059, id_4056, id_4067);
not ( id_6239, id_6233);
nand ( id_6242, id_6233, id_6240);
nand ( id_6253, id_6251, id_6252);
nand ( id_7111, id_7109, id_7110);
nand ( id_7121, id_7119, id_7120);
nand ( id_984, id_5084, id_5087);
nand ( id_987, id_5094, id_5097);
nand ( id_1775, id_5654, id_5657);
nand ( id_1778, id_5664, id_5667);
not ( id_5743, id_5737);
nand ( id_6241, id_6236, id_6239);
or ( id_6329, id_2844, id_2845, id_2846, id_2847);
or ( id_7197, id_4083, id_4084, id_4085, id_4086);
nand ( id_986, id_984, id_985);
nand ( id_989, id_987, id_988);
nand ( id_1777, id_1775, id_1776);
nand ( id_1780, id_1778, id_1779);
not ( id_6259, id_6253);
nand ( id_2841, id_6253, id_6260);
not ( id_7117, id_7111);
nand ( id_4077, id_7111, id_7118);
not ( id_7127, id_7121);
nand ( id_4080, id_7121, id_7128);
nand ( id_6243, id_6241, id_6242);
not ( id_990, id_989);
and ( id_996, id_975, id_986);
not ( id_1781, id_1780);
and ( id_1787, id_1766, id_1777);
nand ( id_2840, id_6256, id_6259);
not ( id_6335, id_6329);
nand ( id_4076, id_7114, id_7117);
nand ( id_4079, id_7124, id_7127);
not ( id_7203, id_7197);
and ( id_995, id_990, id_980);
and ( id_1786, id_1781, id_1771);
not ( id_6249, id_6243);
nand ( id_2838, id_6243, id_6250);
nand ( id_2842, id_2840, id_2841);
nand ( id_4078, id_4076, id_4077);
nand ( id_4081, id_4079, id_4080);
nand ( id_2837, id_6246, id_6249);
not ( id_2843, id_2842);
not ( id_4082, id_4081);
and ( id_4088, id_4067, id_4078);
or ( id_5170, id_995, id_996);
or ( id_5740, id_1786, id_1787);
nand ( id_2839, id_2837, id_2838);
and ( id_2848, id_2843, id_2833);
and ( id_4087, id_4082, id_4072);
nand ( id_1791, id_5740, id_5743);
nand ( id_1003, id_5170, id_5173);
not ( id_5174, id_5170);
not ( id_5744, id_5740);
and ( id_2849, id_2828, id_2839);
or ( id_7200, id_4087, id_4088);
nand ( id_1792, id_5737, id_5744);
nand ( id_1004, id_5167, id_5174);
or ( id_6332, id_2848, id_2849);
nand ( id_320, id_1791, id_1792);
nand ( id_337, id_1003, id_1004);
nand ( id_4092, id_7200, id_7203);
not ( id_7204, id_7200);
not ( id_321, id_320);
not ( id_338, id_337);
nand ( id_4093, id_7197, id_7204);
nand ( id_2855, id_6332, id_6335);
not ( id_6336, id_6332);
nand ( id_369, id_4092, id_4093);
nand ( id_2856, id_6329, id_6336);
not ( id_370, id_369);
nand ( id_398, id_2855, id_2856);
not ( id_399, id_398);

endmodule
